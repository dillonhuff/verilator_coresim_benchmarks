

module coreir_and #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 & in1;

endmodule //coreir_and

module coreir_reg #(parameter init=1, parameter width=1) (
  input clk,
  input [width-1:0] in,
  output [width-1:0] out
);
reg [width-1:0] outReg=init;
always @(posedge clk) begin
  outReg <= in;
end
assign out = outReg;

endmodule //coreir_reg

module coreir_or #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output [width-1:0] out
);
  assign out = in0 | in1;

endmodule //coreir_or

module manyOps (
  input  clk,
  input [15:0] in_0,
  input [15:0] in_1,
  input [15:0] in_10,
  input [15:0] in_100,
  input [15:0] in_1000,
  input [15:0] in_1001,
  input [15:0] in_1002,
  input [15:0] in_1003,
  input [15:0] in_1004,
  input [15:0] in_1005,
  input [15:0] in_1006,
  input [15:0] in_1007,
  input [15:0] in_1008,
  input [15:0] in_1009,
  input [15:0] in_101,
  input [15:0] in_1010,
  input [15:0] in_1011,
  input [15:0] in_1012,
  input [15:0] in_1013,
  input [15:0] in_1014,
  input [15:0] in_1015,
  input [15:0] in_1016,
  input [15:0] in_1017,
  input [15:0] in_1018,
  input [15:0] in_1019,
  input [15:0] in_102,
  input [15:0] in_1020,
  input [15:0] in_1021,
  input [15:0] in_1022,
  input [15:0] in_1023,
  input [15:0] in_1024,
  input [15:0] in_1025,
  input [15:0] in_1026,
  input [15:0] in_1027,
  input [15:0] in_1028,
  input [15:0] in_1029,
  input [15:0] in_103,
  input [15:0] in_1030,
  input [15:0] in_1031,
  input [15:0] in_1032,
  input [15:0] in_1033,
  input [15:0] in_1034,
  input [15:0] in_1035,
  input [15:0] in_1036,
  input [15:0] in_1037,
  input [15:0] in_1038,
  input [15:0] in_1039,
  input [15:0] in_104,
  input [15:0] in_1040,
  input [15:0] in_1041,
  input [15:0] in_1042,
  input [15:0] in_1043,
  input [15:0] in_1044,
  input [15:0] in_1045,
  input [15:0] in_1046,
  input [15:0] in_1047,
  input [15:0] in_1048,
  input [15:0] in_1049,
  input [15:0] in_105,
  input [15:0] in_1050,
  input [15:0] in_1051,
  input [15:0] in_1052,
  input [15:0] in_1053,
  input [15:0] in_1054,
  input [15:0] in_1055,
  input [15:0] in_1056,
  input [15:0] in_1057,
  input [15:0] in_1058,
  input [15:0] in_1059,
  input [15:0] in_106,
  input [15:0] in_1060,
  input [15:0] in_1061,
  input [15:0] in_1062,
  input [15:0] in_1063,
  input [15:0] in_1064,
  input [15:0] in_1065,
  input [15:0] in_1066,
  input [15:0] in_1067,
  input [15:0] in_1068,
  input [15:0] in_1069,
  input [15:0] in_107,
  input [15:0] in_1070,
  input [15:0] in_1071,
  input [15:0] in_1072,
  input [15:0] in_1073,
  input [15:0] in_1074,
  input [15:0] in_1075,
  input [15:0] in_1076,
  input [15:0] in_1077,
  input [15:0] in_1078,
  input [15:0] in_1079,
  input [15:0] in_108,
  input [15:0] in_1080,
  input [15:0] in_1081,
  input [15:0] in_1082,
  input [15:0] in_1083,
  input [15:0] in_1084,
  input [15:0] in_1085,
  input [15:0] in_1086,
  input [15:0] in_1087,
  input [15:0] in_1088,
  input [15:0] in_1089,
  input [15:0] in_109,
  input [15:0] in_1090,
  input [15:0] in_1091,
  input [15:0] in_1092,
  input [15:0] in_1093,
  input [15:0] in_1094,
  input [15:0] in_1095,
  input [15:0] in_1096,
  input [15:0] in_1097,
  input [15:0] in_1098,
  input [15:0] in_1099,
  input [15:0] in_11,
  input [15:0] in_110,
  input [15:0] in_1100,
  input [15:0] in_1101,
  input [15:0] in_1102,
  input [15:0] in_1103,
  input [15:0] in_1104,
  input [15:0] in_1105,
  input [15:0] in_1106,
  input [15:0] in_1107,
  input [15:0] in_1108,
  input [15:0] in_1109,
  input [15:0] in_111,
  input [15:0] in_1110,
  input [15:0] in_1111,
  input [15:0] in_1112,
  input [15:0] in_1113,
  input [15:0] in_1114,
  input [15:0] in_1115,
  input [15:0] in_1116,
  input [15:0] in_1117,
  input [15:0] in_1118,
  input [15:0] in_1119,
  input [15:0] in_112,
  input [15:0] in_1120,
  input [15:0] in_1121,
  input [15:0] in_1122,
  input [15:0] in_1123,
  input [15:0] in_1124,
  input [15:0] in_1125,
  input [15:0] in_1126,
  input [15:0] in_1127,
  input [15:0] in_1128,
  input [15:0] in_1129,
  input [15:0] in_113,
  input [15:0] in_1130,
  input [15:0] in_1131,
  input [15:0] in_1132,
  input [15:0] in_1133,
  input [15:0] in_1134,
  input [15:0] in_1135,
  input [15:0] in_1136,
  input [15:0] in_1137,
  input [15:0] in_1138,
  input [15:0] in_1139,
  input [15:0] in_114,
  input [15:0] in_1140,
  input [15:0] in_1141,
  input [15:0] in_1142,
  input [15:0] in_1143,
  input [15:0] in_1144,
  input [15:0] in_1145,
  input [15:0] in_1146,
  input [15:0] in_1147,
  input [15:0] in_1148,
  input [15:0] in_1149,
  input [15:0] in_115,
  input [15:0] in_1150,
  input [15:0] in_1151,
  input [15:0] in_1152,
  input [15:0] in_1153,
  input [15:0] in_1154,
  input [15:0] in_1155,
  input [15:0] in_1156,
  input [15:0] in_1157,
  input [15:0] in_1158,
  input [15:0] in_1159,
  input [15:0] in_116,
  input [15:0] in_1160,
  input [15:0] in_1161,
  input [15:0] in_1162,
  input [15:0] in_1163,
  input [15:0] in_1164,
  input [15:0] in_1165,
  input [15:0] in_1166,
  input [15:0] in_1167,
  input [15:0] in_1168,
  input [15:0] in_1169,
  input [15:0] in_117,
  input [15:0] in_1170,
  input [15:0] in_1171,
  input [15:0] in_1172,
  input [15:0] in_1173,
  input [15:0] in_1174,
  input [15:0] in_1175,
  input [15:0] in_1176,
  input [15:0] in_1177,
  input [15:0] in_1178,
  input [15:0] in_1179,
  input [15:0] in_118,
  input [15:0] in_1180,
  input [15:0] in_1181,
  input [15:0] in_1182,
  input [15:0] in_1183,
  input [15:0] in_1184,
  input [15:0] in_1185,
  input [15:0] in_1186,
  input [15:0] in_1187,
  input [15:0] in_1188,
  input [15:0] in_1189,
  input [15:0] in_119,
  input [15:0] in_1190,
  input [15:0] in_1191,
  input [15:0] in_1192,
  input [15:0] in_1193,
  input [15:0] in_1194,
  input [15:0] in_1195,
  input [15:0] in_1196,
  input [15:0] in_1197,
  input [15:0] in_1198,
  input [15:0] in_1199,
  input [15:0] in_12,
  input [15:0] in_120,
  input [15:0] in_1200,
  input [15:0] in_1201,
  input [15:0] in_1202,
  input [15:0] in_1203,
  input [15:0] in_1204,
  input [15:0] in_1205,
  input [15:0] in_1206,
  input [15:0] in_1207,
  input [15:0] in_1208,
  input [15:0] in_1209,
  input [15:0] in_121,
  input [15:0] in_1210,
  input [15:0] in_1211,
  input [15:0] in_1212,
  input [15:0] in_1213,
  input [15:0] in_1214,
  input [15:0] in_1215,
  input [15:0] in_1216,
  input [15:0] in_1217,
  input [15:0] in_1218,
  input [15:0] in_1219,
  input [15:0] in_122,
  input [15:0] in_1220,
  input [15:0] in_1221,
  input [15:0] in_1222,
  input [15:0] in_1223,
  input [15:0] in_1224,
  input [15:0] in_1225,
  input [15:0] in_1226,
  input [15:0] in_1227,
  input [15:0] in_1228,
  input [15:0] in_1229,
  input [15:0] in_123,
  input [15:0] in_1230,
  input [15:0] in_1231,
  input [15:0] in_1232,
  input [15:0] in_1233,
  input [15:0] in_1234,
  input [15:0] in_1235,
  input [15:0] in_1236,
  input [15:0] in_1237,
  input [15:0] in_1238,
  input [15:0] in_1239,
  input [15:0] in_124,
  input [15:0] in_1240,
  input [15:0] in_1241,
  input [15:0] in_1242,
  input [15:0] in_1243,
  input [15:0] in_1244,
  input [15:0] in_1245,
  input [15:0] in_1246,
  input [15:0] in_1247,
  input [15:0] in_1248,
  input [15:0] in_1249,
  input [15:0] in_125,
  input [15:0] in_1250,
  input [15:0] in_1251,
  input [15:0] in_1252,
  input [15:0] in_1253,
  input [15:0] in_1254,
  input [15:0] in_1255,
  input [15:0] in_1256,
  input [15:0] in_1257,
  input [15:0] in_1258,
  input [15:0] in_1259,
  input [15:0] in_126,
  input [15:0] in_1260,
  input [15:0] in_1261,
  input [15:0] in_1262,
  input [15:0] in_1263,
  input [15:0] in_1264,
  input [15:0] in_1265,
  input [15:0] in_1266,
  input [15:0] in_1267,
  input [15:0] in_1268,
  input [15:0] in_1269,
  input [15:0] in_127,
  input [15:0] in_1270,
  input [15:0] in_1271,
  input [15:0] in_1272,
  input [15:0] in_1273,
  input [15:0] in_1274,
  input [15:0] in_1275,
  input [15:0] in_1276,
  input [15:0] in_1277,
  input [15:0] in_1278,
  input [15:0] in_1279,
  input [15:0] in_128,
  input [15:0] in_1280,
  input [15:0] in_1281,
  input [15:0] in_1282,
  input [15:0] in_1283,
  input [15:0] in_1284,
  input [15:0] in_1285,
  input [15:0] in_1286,
  input [15:0] in_1287,
  input [15:0] in_1288,
  input [15:0] in_1289,
  input [15:0] in_129,
  input [15:0] in_1290,
  input [15:0] in_1291,
  input [15:0] in_1292,
  input [15:0] in_1293,
  input [15:0] in_1294,
  input [15:0] in_1295,
  input [15:0] in_1296,
  input [15:0] in_1297,
  input [15:0] in_1298,
  input [15:0] in_1299,
  input [15:0] in_13,
  input [15:0] in_130,
  input [15:0] in_1300,
  input [15:0] in_1301,
  input [15:0] in_1302,
  input [15:0] in_1303,
  input [15:0] in_1304,
  input [15:0] in_1305,
  input [15:0] in_1306,
  input [15:0] in_1307,
  input [15:0] in_1308,
  input [15:0] in_1309,
  input [15:0] in_131,
  input [15:0] in_1310,
  input [15:0] in_1311,
  input [15:0] in_1312,
  input [15:0] in_1313,
  input [15:0] in_1314,
  input [15:0] in_1315,
  input [15:0] in_1316,
  input [15:0] in_1317,
  input [15:0] in_1318,
  input [15:0] in_1319,
  input [15:0] in_132,
  input [15:0] in_1320,
  input [15:0] in_1321,
  input [15:0] in_1322,
  input [15:0] in_1323,
  input [15:0] in_1324,
  input [15:0] in_1325,
  input [15:0] in_1326,
  input [15:0] in_1327,
  input [15:0] in_1328,
  input [15:0] in_1329,
  input [15:0] in_133,
  input [15:0] in_1330,
  input [15:0] in_1331,
  input [15:0] in_1332,
  input [15:0] in_1333,
  input [15:0] in_1334,
  input [15:0] in_1335,
  input [15:0] in_1336,
  input [15:0] in_1337,
  input [15:0] in_1338,
  input [15:0] in_1339,
  input [15:0] in_134,
  input [15:0] in_1340,
  input [15:0] in_1341,
  input [15:0] in_1342,
  input [15:0] in_1343,
  input [15:0] in_1344,
  input [15:0] in_1345,
  input [15:0] in_1346,
  input [15:0] in_1347,
  input [15:0] in_1348,
  input [15:0] in_1349,
  input [15:0] in_135,
  input [15:0] in_1350,
  input [15:0] in_1351,
  input [15:0] in_1352,
  input [15:0] in_1353,
  input [15:0] in_1354,
  input [15:0] in_1355,
  input [15:0] in_1356,
  input [15:0] in_1357,
  input [15:0] in_1358,
  input [15:0] in_1359,
  input [15:0] in_136,
  input [15:0] in_1360,
  input [15:0] in_1361,
  input [15:0] in_1362,
  input [15:0] in_1363,
  input [15:0] in_1364,
  input [15:0] in_1365,
  input [15:0] in_1366,
  input [15:0] in_1367,
  input [15:0] in_1368,
  input [15:0] in_1369,
  input [15:0] in_137,
  input [15:0] in_1370,
  input [15:0] in_1371,
  input [15:0] in_1372,
  input [15:0] in_1373,
  input [15:0] in_1374,
  input [15:0] in_1375,
  input [15:0] in_1376,
  input [15:0] in_1377,
  input [15:0] in_1378,
  input [15:0] in_1379,
  input [15:0] in_138,
  input [15:0] in_1380,
  input [15:0] in_1381,
  input [15:0] in_1382,
  input [15:0] in_1383,
  input [15:0] in_1384,
  input [15:0] in_1385,
  input [15:0] in_1386,
  input [15:0] in_1387,
  input [15:0] in_1388,
  input [15:0] in_1389,
  input [15:0] in_139,
  input [15:0] in_1390,
  input [15:0] in_1391,
  input [15:0] in_1392,
  input [15:0] in_1393,
  input [15:0] in_1394,
  input [15:0] in_1395,
  input [15:0] in_1396,
  input [15:0] in_1397,
  input [15:0] in_1398,
  input [15:0] in_1399,
  input [15:0] in_14,
  input [15:0] in_140,
  input [15:0] in_1400,
  input [15:0] in_1401,
  input [15:0] in_1402,
  input [15:0] in_1403,
  input [15:0] in_1404,
  input [15:0] in_1405,
  input [15:0] in_1406,
  input [15:0] in_1407,
  input [15:0] in_1408,
  input [15:0] in_1409,
  input [15:0] in_141,
  input [15:0] in_1410,
  input [15:0] in_1411,
  input [15:0] in_1412,
  input [15:0] in_1413,
  input [15:0] in_1414,
  input [15:0] in_1415,
  input [15:0] in_1416,
  input [15:0] in_1417,
  input [15:0] in_1418,
  input [15:0] in_1419,
  input [15:0] in_142,
  input [15:0] in_1420,
  input [15:0] in_1421,
  input [15:0] in_1422,
  input [15:0] in_1423,
  input [15:0] in_1424,
  input [15:0] in_1425,
  input [15:0] in_1426,
  input [15:0] in_1427,
  input [15:0] in_1428,
  input [15:0] in_1429,
  input [15:0] in_143,
  input [15:0] in_1430,
  input [15:0] in_1431,
  input [15:0] in_1432,
  input [15:0] in_1433,
  input [15:0] in_1434,
  input [15:0] in_1435,
  input [15:0] in_1436,
  input [15:0] in_1437,
  input [15:0] in_1438,
  input [15:0] in_1439,
  input [15:0] in_144,
  input [15:0] in_1440,
  input [15:0] in_1441,
  input [15:0] in_1442,
  input [15:0] in_1443,
  input [15:0] in_1444,
  input [15:0] in_1445,
  input [15:0] in_1446,
  input [15:0] in_1447,
  input [15:0] in_1448,
  input [15:0] in_1449,
  input [15:0] in_145,
  input [15:0] in_1450,
  input [15:0] in_1451,
  input [15:0] in_1452,
  input [15:0] in_1453,
  input [15:0] in_1454,
  input [15:0] in_1455,
  input [15:0] in_1456,
  input [15:0] in_1457,
  input [15:0] in_1458,
  input [15:0] in_1459,
  input [15:0] in_146,
  input [15:0] in_1460,
  input [15:0] in_1461,
  input [15:0] in_1462,
  input [15:0] in_1463,
  input [15:0] in_1464,
  input [15:0] in_1465,
  input [15:0] in_1466,
  input [15:0] in_1467,
  input [15:0] in_1468,
  input [15:0] in_1469,
  input [15:0] in_147,
  input [15:0] in_1470,
  input [15:0] in_1471,
  input [15:0] in_1472,
  input [15:0] in_1473,
  input [15:0] in_1474,
  input [15:0] in_1475,
  input [15:0] in_1476,
  input [15:0] in_1477,
  input [15:0] in_1478,
  input [15:0] in_1479,
  input [15:0] in_148,
  input [15:0] in_1480,
  input [15:0] in_1481,
  input [15:0] in_1482,
  input [15:0] in_1483,
  input [15:0] in_1484,
  input [15:0] in_1485,
  input [15:0] in_1486,
  input [15:0] in_1487,
  input [15:0] in_1488,
  input [15:0] in_1489,
  input [15:0] in_149,
  input [15:0] in_1490,
  input [15:0] in_1491,
  input [15:0] in_1492,
  input [15:0] in_1493,
  input [15:0] in_1494,
  input [15:0] in_1495,
  input [15:0] in_1496,
  input [15:0] in_1497,
  input [15:0] in_1498,
  input [15:0] in_1499,
  input [15:0] in_15,
  input [15:0] in_150,
  input [15:0] in_1500,
  input [15:0] in_1501,
  input [15:0] in_1502,
  input [15:0] in_1503,
  input [15:0] in_1504,
  input [15:0] in_1505,
  input [15:0] in_1506,
  input [15:0] in_1507,
  input [15:0] in_1508,
  input [15:0] in_1509,
  input [15:0] in_151,
  input [15:0] in_1510,
  input [15:0] in_1511,
  input [15:0] in_1512,
  input [15:0] in_1513,
  input [15:0] in_1514,
  input [15:0] in_1515,
  input [15:0] in_1516,
  input [15:0] in_1517,
  input [15:0] in_1518,
  input [15:0] in_1519,
  input [15:0] in_152,
  input [15:0] in_1520,
  input [15:0] in_1521,
  input [15:0] in_1522,
  input [15:0] in_1523,
  input [15:0] in_1524,
  input [15:0] in_1525,
  input [15:0] in_1526,
  input [15:0] in_1527,
  input [15:0] in_1528,
  input [15:0] in_1529,
  input [15:0] in_153,
  input [15:0] in_1530,
  input [15:0] in_1531,
  input [15:0] in_1532,
  input [15:0] in_1533,
  input [15:0] in_1534,
  input [15:0] in_1535,
  input [15:0] in_1536,
  input [15:0] in_1537,
  input [15:0] in_1538,
  input [15:0] in_1539,
  input [15:0] in_154,
  input [15:0] in_1540,
  input [15:0] in_1541,
  input [15:0] in_1542,
  input [15:0] in_1543,
  input [15:0] in_1544,
  input [15:0] in_1545,
  input [15:0] in_1546,
  input [15:0] in_1547,
  input [15:0] in_1548,
  input [15:0] in_1549,
  input [15:0] in_155,
  input [15:0] in_1550,
  input [15:0] in_1551,
  input [15:0] in_1552,
  input [15:0] in_1553,
  input [15:0] in_1554,
  input [15:0] in_1555,
  input [15:0] in_1556,
  input [15:0] in_1557,
  input [15:0] in_1558,
  input [15:0] in_1559,
  input [15:0] in_156,
  input [15:0] in_1560,
  input [15:0] in_1561,
  input [15:0] in_1562,
  input [15:0] in_1563,
  input [15:0] in_1564,
  input [15:0] in_1565,
  input [15:0] in_1566,
  input [15:0] in_1567,
  input [15:0] in_1568,
  input [15:0] in_1569,
  input [15:0] in_157,
  input [15:0] in_1570,
  input [15:0] in_1571,
  input [15:0] in_1572,
  input [15:0] in_1573,
  input [15:0] in_1574,
  input [15:0] in_1575,
  input [15:0] in_1576,
  input [15:0] in_1577,
  input [15:0] in_1578,
  input [15:0] in_1579,
  input [15:0] in_158,
  input [15:0] in_1580,
  input [15:0] in_1581,
  input [15:0] in_1582,
  input [15:0] in_1583,
  input [15:0] in_1584,
  input [15:0] in_1585,
  input [15:0] in_1586,
  input [15:0] in_1587,
  input [15:0] in_1588,
  input [15:0] in_1589,
  input [15:0] in_159,
  input [15:0] in_1590,
  input [15:0] in_1591,
  input [15:0] in_1592,
  input [15:0] in_1593,
  input [15:0] in_1594,
  input [15:0] in_1595,
  input [15:0] in_1596,
  input [15:0] in_1597,
  input [15:0] in_1598,
  input [15:0] in_1599,
  input [15:0] in_16,
  input [15:0] in_160,
  input [15:0] in_1600,
  input [15:0] in_1601,
  input [15:0] in_1602,
  input [15:0] in_1603,
  input [15:0] in_1604,
  input [15:0] in_1605,
  input [15:0] in_1606,
  input [15:0] in_1607,
  input [15:0] in_1608,
  input [15:0] in_1609,
  input [15:0] in_161,
  input [15:0] in_1610,
  input [15:0] in_1611,
  input [15:0] in_1612,
  input [15:0] in_1613,
  input [15:0] in_1614,
  input [15:0] in_1615,
  input [15:0] in_1616,
  input [15:0] in_1617,
  input [15:0] in_1618,
  input [15:0] in_1619,
  input [15:0] in_162,
  input [15:0] in_1620,
  input [15:0] in_1621,
  input [15:0] in_1622,
  input [15:0] in_1623,
  input [15:0] in_1624,
  input [15:0] in_1625,
  input [15:0] in_1626,
  input [15:0] in_1627,
  input [15:0] in_1628,
  input [15:0] in_1629,
  input [15:0] in_163,
  input [15:0] in_1630,
  input [15:0] in_1631,
  input [15:0] in_1632,
  input [15:0] in_1633,
  input [15:0] in_1634,
  input [15:0] in_1635,
  input [15:0] in_1636,
  input [15:0] in_1637,
  input [15:0] in_1638,
  input [15:0] in_1639,
  input [15:0] in_164,
  input [15:0] in_1640,
  input [15:0] in_1641,
  input [15:0] in_1642,
  input [15:0] in_1643,
  input [15:0] in_1644,
  input [15:0] in_1645,
  input [15:0] in_1646,
  input [15:0] in_1647,
  input [15:0] in_1648,
  input [15:0] in_1649,
  input [15:0] in_165,
  input [15:0] in_1650,
  input [15:0] in_1651,
  input [15:0] in_1652,
  input [15:0] in_1653,
  input [15:0] in_1654,
  input [15:0] in_1655,
  input [15:0] in_1656,
  input [15:0] in_1657,
  input [15:0] in_1658,
  input [15:0] in_1659,
  input [15:0] in_166,
  input [15:0] in_1660,
  input [15:0] in_1661,
  input [15:0] in_1662,
  input [15:0] in_1663,
  input [15:0] in_1664,
  input [15:0] in_1665,
  input [15:0] in_1666,
  input [15:0] in_1667,
  input [15:0] in_1668,
  input [15:0] in_1669,
  input [15:0] in_167,
  input [15:0] in_1670,
  input [15:0] in_1671,
  input [15:0] in_1672,
  input [15:0] in_1673,
  input [15:0] in_1674,
  input [15:0] in_1675,
  input [15:0] in_1676,
  input [15:0] in_1677,
  input [15:0] in_1678,
  input [15:0] in_1679,
  input [15:0] in_168,
  input [15:0] in_1680,
  input [15:0] in_1681,
  input [15:0] in_1682,
  input [15:0] in_1683,
  input [15:0] in_1684,
  input [15:0] in_1685,
  input [15:0] in_1686,
  input [15:0] in_1687,
  input [15:0] in_1688,
  input [15:0] in_1689,
  input [15:0] in_169,
  input [15:0] in_1690,
  input [15:0] in_1691,
  input [15:0] in_1692,
  input [15:0] in_1693,
  input [15:0] in_1694,
  input [15:0] in_1695,
  input [15:0] in_1696,
  input [15:0] in_1697,
  input [15:0] in_1698,
  input [15:0] in_1699,
  input [15:0] in_17,
  input [15:0] in_170,
  input [15:0] in_1700,
  input [15:0] in_1701,
  input [15:0] in_1702,
  input [15:0] in_1703,
  input [15:0] in_1704,
  input [15:0] in_1705,
  input [15:0] in_1706,
  input [15:0] in_1707,
  input [15:0] in_1708,
  input [15:0] in_1709,
  input [15:0] in_171,
  input [15:0] in_1710,
  input [15:0] in_1711,
  input [15:0] in_1712,
  input [15:0] in_1713,
  input [15:0] in_1714,
  input [15:0] in_1715,
  input [15:0] in_1716,
  input [15:0] in_1717,
  input [15:0] in_1718,
  input [15:0] in_1719,
  input [15:0] in_172,
  input [15:0] in_1720,
  input [15:0] in_1721,
  input [15:0] in_1722,
  input [15:0] in_1723,
  input [15:0] in_1724,
  input [15:0] in_1725,
  input [15:0] in_1726,
  input [15:0] in_1727,
  input [15:0] in_1728,
  input [15:0] in_1729,
  input [15:0] in_173,
  input [15:0] in_1730,
  input [15:0] in_1731,
  input [15:0] in_1732,
  input [15:0] in_1733,
  input [15:0] in_1734,
  input [15:0] in_1735,
  input [15:0] in_1736,
  input [15:0] in_1737,
  input [15:0] in_1738,
  input [15:0] in_1739,
  input [15:0] in_174,
  input [15:0] in_1740,
  input [15:0] in_1741,
  input [15:0] in_1742,
  input [15:0] in_1743,
  input [15:0] in_1744,
  input [15:0] in_1745,
  input [15:0] in_1746,
  input [15:0] in_1747,
  input [15:0] in_1748,
  input [15:0] in_1749,
  input [15:0] in_175,
  input [15:0] in_1750,
  input [15:0] in_1751,
  input [15:0] in_1752,
  input [15:0] in_1753,
  input [15:0] in_1754,
  input [15:0] in_1755,
  input [15:0] in_1756,
  input [15:0] in_1757,
  input [15:0] in_1758,
  input [15:0] in_1759,
  input [15:0] in_176,
  input [15:0] in_1760,
  input [15:0] in_1761,
  input [15:0] in_1762,
  input [15:0] in_1763,
  input [15:0] in_1764,
  input [15:0] in_1765,
  input [15:0] in_1766,
  input [15:0] in_1767,
  input [15:0] in_1768,
  input [15:0] in_1769,
  input [15:0] in_177,
  input [15:0] in_1770,
  input [15:0] in_1771,
  input [15:0] in_1772,
  input [15:0] in_1773,
  input [15:0] in_1774,
  input [15:0] in_1775,
  input [15:0] in_1776,
  input [15:0] in_1777,
  input [15:0] in_1778,
  input [15:0] in_1779,
  input [15:0] in_178,
  input [15:0] in_1780,
  input [15:0] in_1781,
  input [15:0] in_1782,
  input [15:0] in_1783,
  input [15:0] in_1784,
  input [15:0] in_1785,
  input [15:0] in_1786,
  input [15:0] in_1787,
  input [15:0] in_1788,
  input [15:0] in_1789,
  input [15:0] in_179,
  input [15:0] in_1790,
  input [15:0] in_1791,
  input [15:0] in_1792,
  input [15:0] in_1793,
  input [15:0] in_1794,
  input [15:0] in_1795,
  input [15:0] in_1796,
  input [15:0] in_1797,
  input [15:0] in_1798,
  input [15:0] in_1799,
  input [15:0] in_18,
  input [15:0] in_180,
  input [15:0] in_1800,
  input [15:0] in_1801,
  input [15:0] in_1802,
  input [15:0] in_1803,
  input [15:0] in_1804,
  input [15:0] in_1805,
  input [15:0] in_1806,
  input [15:0] in_1807,
  input [15:0] in_1808,
  input [15:0] in_1809,
  input [15:0] in_181,
  input [15:0] in_1810,
  input [15:0] in_1811,
  input [15:0] in_1812,
  input [15:0] in_1813,
  input [15:0] in_1814,
  input [15:0] in_1815,
  input [15:0] in_1816,
  input [15:0] in_1817,
  input [15:0] in_1818,
  input [15:0] in_1819,
  input [15:0] in_182,
  input [15:0] in_1820,
  input [15:0] in_1821,
  input [15:0] in_1822,
  input [15:0] in_1823,
  input [15:0] in_1824,
  input [15:0] in_1825,
  input [15:0] in_1826,
  input [15:0] in_1827,
  input [15:0] in_1828,
  input [15:0] in_1829,
  input [15:0] in_183,
  input [15:0] in_1830,
  input [15:0] in_1831,
  input [15:0] in_1832,
  input [15:0] in_1833,
  input [15:0] in_1834,
  input [15:0] in_1835,
  input [15:0] in_1836,
  input [15:0] in_1837,
  input [15:0] in_1838,
  input [15:0] in_1839,
  input [15:0] in_184,
  input [15:0] in_1840,
  input [15:0] in_1841,
  input [15:0] in_1842,
  input [15:0] in_1843,
  input [15:0] in_1844,
  input [15:0] in_1845,
  input [15:0] in_1846,
  input [15:0] in_1847,
  input [15:0] in_1848,
  input [15:0] in_1849,
  input [15:0] in_185,
  input [15:0] in_1850,
  input [15:0] in_1851,
  input [15:0] in_1852,
  input [15:0] in_1853,
  input [15:0] in_1854,
  input [15:0] in_1855,
  input [15:0] in_1856,
  input [15:0] in_1857,
  input [15:0] in_1858,
  input [15:0] in_1859,
  input [15:0] in_186,
  input [15:0] in_1860,
  input [15:0] in_1861,
  input [15:0] in_1862,
  input [15:0] in_1863,
  input [15:0] in_1864,
  input [15:0] in_1865,
  input [15:0] in_1866,
  input [15:0] in_1867,
  input [15:0] in_1868,
  input [15:0] in_1869,
  input [15:0] in_187,
  input [15:0] in_1870,
  input [15:0] in_1871,
  input [15:0] in_1872,
  input [15:0] in_1873,
  input [15:0] in_1874,
  input [15:0] in_1875,
  input [15:0] in_1876,
  input [15:0] in_1877,
  input [15:0] in_1878,
  input [15:0] in_1879,
  input [15:0] in_188,
  input [15:0] in_1880,
  input [15:0] in_1881,
  input [15:0] in_1882,
  input [15:0] in_1883,
  input [15:0] in_1884,
  input [15:0] in_1885,
  input [15:0] in_1886,
  input [15:0] in_1887,
  input [15:0] in_1888,
  input [15:0] in_1889,
  input [15:0] in_189,
  input [15:0] in_1890,
  input [15:0] in_1891,
  input [15:0] in_1892,
  input [15:0] in_1893,
  input [15:0] in_1894,
  input [15:0] in_1895,
  input [15:0] in_1896,
  input [15:0] in_1897,
  input [15:0] in_1898,
  input [15:0] in_1899,
  input [15:0] in_19,
  input [15:0] in_190,
  input [15:0] in_1900,
  input [15:0] in_1901,
  input [15:0] in_1902,
  input [15:0] in_1903,
  input [15:0] in_1904,
  input [15:0] in_1905,
  input [15:0] in_1906,
  input [15:0] in_1907,
  input [15:0] in_1908,
  input [15:0] in_1909,
  input [15:0] in_191,
  input [15:0] in_1910,
  input [15:0] in_1911,
  input [15:0] in_1912,
  input [15:0] in_1913,
  input [15:0] in_1914,
  input [15:0] in_1915,
  input [15:0] in_1916,
  input [15:0] in_1917,
  input [15:0] in_1918,
  input [15:0] in_1919,
  input [15:0] in_192,
  input [15:0] in_1920,
  input [15:0] in_1921,
  input [15:0] in_1922,
  input [15:0] in_1923,
  input [15:0] in_1924,
  input [15:0] in_1925,
  input [15:0] in_1926,
  input [15:0] in_1927,
  input [15:0] in_1928,
  input [15:0] in_1929,
  input [15:0] in_193,
  input [15:0] in_1930,
  input [15:0] in_1931,
  input [15:0] in_1932,
  input [15:0] in_1933,
  input [15:0] in_1934,
  input [15:0] in_1935,
  input [15:0] in_1936,
  input [15:0] in_1937,
  input [15:0] in_1938,
  input [15:0] in_1939,
  input [15:0] in_194,
  input [15:0] in_1940,
  input [15:0] in_1941,
  input [15:0] in_1942,
  input [15:0] in_1943,
  input [15:0] in_1944,
  input [15:0] in_1945,
  input [15:0] in_1946,
  input [15:0] in_1947,
  input [15:0] in_1948,
  input [15:0] in_1949,
  input [15:0] in_195,
  input [15:0] in_1950,
  input [15:0] in_1951,
  input [15:0] in_1952,
  input [15:0] in_1953,
  input [15:0] in_1954,
  input [15:0] in_1955,
  input [15:0] in_1956,
  input [15:0] in_1957,
  input [15:0] in_1958,
  input [15:0] in_1959,
  input [15:0] in_196,
  input [15:0] in_1960,
  input [15:0] in_1961,
  input [15:0] in_1962,
  input [15:0] in_1963,
  input [15:0] in_1964,
  input [15:0] in_1965,
  input [15:0] in_1966,
  input [15:0] in_1967,
  input [15:0] in_1968,
  input [15:0] in_1969,
  input [15:0] in_197,
  input [15:0] in_1970,
  input [15:0] in_1971,
  input [15:0] in_1972,
  input [15:0] in_1973,
  input [15:0] in_1974,
  input [15:0] in_1975,
  input [15:0] in_1976,
  input [15:0] in_1977,
  input [15:0] in_1978,
  input [15:0] in_1979,
  input [15:0] in_198,
  input [15:0] in_1980,
  input [15:0] in_1981,
  input [15:0] in_1982,
  input [15:0] in_1983,
  input [15:0] in_1984,
  input [15:0] in_1985,
  input [15:0] in_1986,
  input [15:0] in_1987,
  input [15:0] in_1988,
  input [15:0] in_1989,
  input [15:0] in_199,
  input [15:0] in_1990,
  input [15:0] in_1991,
  input [15:0] in_1992,
  input [15:0] in_1993,
  input [15:0] in_1994,
  input [15:0] in_1995,
  input [15:0] in_1996,
  input [15:0] in_1997,
  input [15:0] in_1998,
  input [15:0] in_1999,
  input [15:0] in_2,
  input [15:0] in_20,
  input [15:0] in_200,
  input [15:0] in_201,
  input [15:0] in_202,
  input [15:0] in_203,
  input [15:0] in_204,
  input [15:0] in_205,
  input [15:0] in_206,
  input [15:0] in_207,
  input [15:0] in_208,
  input [15:0] in_209,
  input [15:0] in_21,
  input [15:0] in_210,
  input [15:0] in_211,
  input [15:0] in_212,
  input [15:0] in_213,
  input [15:0] in_214,
  input [15:0] in_215,
  input [15:0] in_216,
  input [15:0] in_217,
  input [15:0] in_218,
  input [15:0] in_219,
  input [15:0] in_22,
  input [15:0] in_220,
  input [15:0] in_221,
  input [15:0] in_222,
  input [15:0] in_223,
  input [15:0] in_224,
  input [15:0] in_225,
  input [15:0] in_226,
  input [15:0] in_227,
  input [15:0] in_228,
  input [15:0] in_229,
  input [15:0] in_23,
  input [15:0] in_230,
  input [15:0] in_231,
  input [15:0] in_232,
  input [15:0] in_233,
  input [15:0] in_234,
  input [15:0] in_235,
  input [15:0] in_236,
  input [15:0] in_237,
  input [15:0] in_238,
  input [15:0] in_239,
  input [15:0] in_24,
  input [15:0] in_240,
  input [15:0] in_241,
  input [15:0] in_242,
  input [15:0] in_243,
  input [15:0] in_244,
  input [15:0] in_245,
  input [15:0] in_246,
  input [15:0] in_247,
  input [15:0] in_248,
  input [15:0] in_249,
  input [15:0] in_25,
  input [15:0] in_250,
  input [15:0] in_251,
  input [15:0] in_252,
  input [15:0] in_253,
  input [15:0] in_254,
  input [15:0] in_255,
  input [15:0] in_256,
  input [15:0] in_257,
  input [15:0] in_258,
  input [15:0] in_259,
  input [15:0] in_26,
  input [15:0] in_260,
  input [15:0] in_261,
  input [15:0] in_262,
  input [15:0] in_263,
  input [15:0] in_264,
  input [15:0] in_265,
  input [15:0] in_266,
  input [15:0] in_267,
  input [15:0] in_268,
  input [15:0] in_269,
  input [15:0] in_27,
  input [15:0] in_270,
  input [15:0] in_271,
  input [15:0] in_272,
  input [15:0] in_273,
  input [15:0] in_274,
  input [15:0] in_275,
  input [15:0] in_276,
  input [15:0] in_277,
  input [15:0] in_278,
  input [15:0] in_279,
  input [15:0] in_28,
  input [15:0] in_280,
  input [15:0] in_281,
  input [15:0] in_282,
  input [15:0] in_283,
  input [15:0] in_284,
  input [15:0] in_285,
  input [15:0] in_286,
  input [15:0] in_287,
  input [15:0] in_288,
  input [15:0] in_289,
  input [15:0] in_29,
  input [15:0] in_290,
  input [15:0] in_291,
  input [15:0] in_292,
  input [15:0] in_293,
  input [15:0] in_294,
  input [15:0] in_295,
  input [15:0] in_296,
  input [15:0] in_297,
  input [15:0] in_298,
  input [15:0] in_299,
  input [15:0] in_3,
  input [15:0] in_30,
  input [15:0] in_300,
  input [15:0] in_301,
  input [15:0] in_302,
  input [15:0] in_303,
  input [15:0] in_304,
  input [15:0] in_305,
  input [15:0] in_306,
  input [15:0] in_307,
  input [15:0] in_308,
  input [15:0] in_309,
  input [15:0] in_31,
  input [15:0] in_310,
  input [15:0] in_311,
  input [15:0] in_312,
  input [15:0] in_313,
  input [15:0] in_314,
  input [15:0] in_315,
  input [15:0] in_316,
  input [15:0] in_317,
  input [15:0] in_318,
  input [15:0] in_319,
  input [15:0] in_32,
  input [15:0] in_320,
  input [15:0] in_321,
  input [15:0] in_322,
  input [15:0] in_323,
  input [15:0] in_324,
  input [15:0] in_325,
  input [15:0] in_326,
  input [15:0] in_327,
  input [15:0] in_328,
  input [15:0] in_329,
  input [15:0] in_33,
  input [15:0] in_330,
  input [15:0] in_331,
  input [15:0] in_332,
  input [15:0] in_333,
  input [15:0] in_334,
  input [15:0] in_335,
  input [15:0] in_336,
  input [15:0] in_337,
  input [15:0] in_338,
  input [15:0] in_339,
  input [15:0] in_34,
  input [15:0] in_340,
  input [15:0] in_341,
  input [15:0] in_342,
  input [15:0] in_343,
  input [15:0] in_344,
  input [15:0] in_345,
  input [15:0] in_346,
  input [15:0] in_347,
  input [15:0] in_348,
  input [15:0] in_349,
  input [15:0] in_35,
  input [15:0] in_350,
  input [15:0] in_351,
  input [15:0] in_352,
  input [15:0] in_353,
  input [15:0] in_354,
  input [15:0] in_355,
  input [15:0] in_356,
  input [15:0] in_357,
  input [15:0] in_358,
  input [15:0] in_359,
  input [15:0] in_36,
  input [15:0] in_360,
  input [15:0] in_361,
  input [15:0] in_362,
  input [15:0] in_363,
  input [15:0] in_364,
  input [15:0] in_365,
  input [15:0] in_366,
  input [15:0] in_367,
  input [15:0] in_368,
  input [15:0] in_369,
  input [15:0] in_37,
  input [15:0] in_370,
  input [15:0] in_371,
  input [15:0] in_372,
  input [15:0] in_373,
  input [15:0] in_374,
  input [15:0] in_375,
  input [15:0] in_376,
  input [15:0] in_377,
  input [15:0] in_378,
  input [15:0] in_379,
  input [15:0] in_38,
  input [15:0] in_380,
  input [15:0] in_381,
  input [15:0] in_382,
  input [15:0] in_383,
  input [15:0] in_384,
  input [15:0] in_385,
  input [15:0] in_386,
  input [15:0] in_387,
  input [15:0] in_388,
  input [15:0] in_389,
  input [15:0] in_39,
  input [15:0] in_390,
  input [15:0] in_391,
  input [15:0] in_392,
  input [15:0] in_393,
  input [15:0] in_394,
  input [15:0] in_395,
  input [15:0] in_396,
  input [15:0] in_397,
  input [15:0] in_398,
  input [15:0] in_399,
  input [15:0] in_4,
  input [15:0] in_40,
  input [15:0] in_400,
  input [15:0] in_401,
  input [15:0] in_402,
  input [15:0] in_403,
  input [15:0] in_404,
  input [15:0] in_405,
  input [15:0] in_406,
  input [15:0] in_407,
  input [15:0] in_408,
  input [15:0] in_409,
  input [15:0] in_41,
  input [15:0] in_410,
  input [15:0] in_411,
  input [15:0] in_412,
  input [15:0] in_413,
  input [15:0] in_414,
  input [15:0] in_415,
  input [15:0] in_416,
  input [15:0] in_417,
  input [15:0] in_418,
  input [15:0] in_419,
  input [15:0] in_42,
  input [15:0] in_420,
  input [15:0] in_421,
  input [15:0] in_422,
  input [15:0] in_423,
  input [15:0] in_424,
  input [15:0] in_425,
  input [15:0] in_426,
  input [15:0] in_427,
  input [15:0] in_428,
  input [15:0] in_429,
  input [15:0] in_43,
  input [15:0] in_430,
  input [15:0] in_431,
  input [15:0] in_432,
  input [15:0] in_433,
  input [15:0] in_434,
  input [15:0] in_435,
  input [15:0] in_436,
  input [15:0] in_437,
  input [15:0] in_438,
  input [15:0] in_439,
  input [15:0] in_44,
  input [15:0] in_440,
  input [15:0] in_441,
  input [15:0] in_442,
  input [15:0] in_443,
  input [15:0] in_444,
  input [15:0] in_445,
  input [15:0] in_446,
  input [15:0] in_447,
  input [15:0] in_448,
  input [15:0] in_449,
  input [15:0] in_45,
  input [15:0] in_450,
  input [15:0] in_451,
  input [15:0] in_452,
  input [15:0] in_453,
  input [15:0] in_454,
  input [15:0] in_455,
  input [15:0] in_456,
  input [15:0] in_457,
  input [15:0] in_458,
  input [15:0] in_459,
  input [15:0] in_46,
  input [15:0] in_460,
  input [15:0] in_461,
  input [15:0] in_462,
  input [15:0] in_463,
  input [15:0] in_464,
  input [15:0] in_465,
  input [15:0] in_466,
  input [15:0] in_467,
  input [15:0] in_468,
  input [15:0] in_469,
  input [15:0] in_47,
  input [15:0] in_470,
  input [15:0] in_471,
  input [15:0] in_472,
  input [15:0] in_473,
  input [15:0] in_474,
  input [15:0] in_475,
  input [15:0] in_476,
  input [15:0] in_477,
  input [15:0] in_478,
  input [15:0] in_479,
  input [15:0] in_48,
  input [15:0] in_480,
  input [15:0] in_481,
  input [15:0] in_482,
  input [15:0] in_483,
  input [15:0] in_484,
  input [15:0] in_485,
  input [15:0] in_486,
  input [15:0] in_487,
  input [15:0] in_488,
  input [15:0] in_489,
  input [15:0] in_49,
  input [15:0] in_490,
  input [15:0] in_491,
  input [15:0] in_492,
  input [15:0] in_493,
  input [15:0] in_494,
  input [15:0] in_495,
  input [15:0] in_496,
  input [15:0] in_497,
  input [15:0] in_498,
  input [15:0] in_499,
  input [15:0] in_5,
  input [15:0] in_50,
  input [15:0] in_500,
  input [15:0] in_501,
  input [15:0] in_502,
  input [15:0] in_503,
  input [15:0] in_504,
  input [15:0] in_505,
  input [15:0] in_506,
  input [15:0] in_507,
  input [15:0] in_508,
  input [15:0] in_509,
  input [15:0] in_51,
  input [15:0] in_510,
  input [15:0] in_511,
  input [15:0] in_512,
  input [15:0] in_513,
  input [15:0] in_514,
  input [15:0] in_515,
  input [15:0] in_516,
  input [15:0] in_517,
  input [15:0] in_518,
  input [15:0] in_519,
  input [15:0] in_52,
  input [15:0] in_520,
  input [15:0] in_521,
  input [15:0] in_522,
  input [15:0] in_523,
  input [15:0] in_524,
  input [15:0] in_525,
  input [15:0] in_526,
  input [15:0] in_527,
  input [15:0] in_528,
  input [15:0] in_529,
  input [15:0] in_53,
  input [15:0] in_530,
  input [15:0] in_531,
  input [15:0] in_532,
  input [15:0] in_533,
  input [15:0] in_534,
  input [15:0] in_535,
  input [15:0] in_536,
  input [15:0] in_537,
  input [15:0] in_538,
  input [15:0] in_539,
  input [15:0] in_54,
  input [15:0] in_540,
  input [15:0] in_541,
  input [15:0] in_542,
  input [15:0] in_543,
  input [15:0] in_544,
  input [15:0] in_545,
  input [15:0] in_546,
  input [15:0] in_547,
  input [15:0] in_548,
  input [15:0] in_549,
  input [15:0] in_55,
  input [15:0] in_550,
  input [15:0] in_551,
  input [15:0] in_552,
  input [15:0] in_553,
  input [15:0] in_554,
  input [15:0] in_555,
  input [15:0] in_556,
  input [15:0] in_557,
  input [15:0] in_558,
  input [15:0] in_559,
  input [15:0] in_56,
  input [15:0] in_560,
  input [15:0] in_561,
  input [15:0] in_562,
  input [15:0] in_563,
  input [15:0] in_564,
  input [15:0] in_565,
  input [15:0] in_566,
  input [15:0] in_567,
  input [15:0] in_568,
  input [15:0] in_569,
  input [15:0] in_57,
  input [15:0] in_570,
  input [15:0] in_571,
  input [15:0] in_572,
  input [15:0] in_573,
  input [15:0] in_574,
  input [15:0] in_575,
  input [15:0] in_576,
  input [15:0] in_577,
  input [15:0] in_578,
  input [15:0] in_579,
  input [15:0] in_58,
  input [15:0] in_580,
  input [15:0] in_581,
  input [15:0] in_582,
  input [15:0] in_583,
  input [15:0] in_584,
  input [15:0] in_585,
  input [15:0] in_586,
  input [15:0] in_587,
  input [15:0] in_588,
  input [15:0] in_589,
  input [15:0] in_59,
  input [15:0] in_590,
  input [15:0] in_591,
  input [15:0] in_592,
  input [15:0] in_593,
  input [15:0] in_594,
  input [15:0] in_595,
  input [15:0] in_596,
  input [15:0] in_597,
  input [15:0] in_598,
  input [15:0] in_599,
  input [15:0] in_6,
  input [15:0] in_60,
  input [15:0] in_600,
  input [15:0] in_601,
  input [15:0] in_602,
  input [15:0] in_603,
  input [15:0] in_604,
  input [15:0] in_605,
  input [15:0] in_606,
  input [15:0] in_607,
  input [15:0] in_608,
  input [15:0] in_609,
  input [15:0] in_61,
  input [15:0] in_610,
  input [15:0] in_611,
  input [15:0] in_612,
  input [15:0] in_613,
  input [15:0] in_614,
  input [15:0] in_615,
  input [15:0] in_616,
  input [15:0] in_617,
  input [15:0] in_618,
  input [15:0] in_619,
  input [15:0] in_62,
  input [15:0] in_620,
  input [15:0] in_621,
  input [15:0] in_622,
  input [15:0] in_623,
  input [15:0] in_624,
  input [15:0] in_625,
  input [15:0] in_626,
  input [15:0] in_627,
  input [15:0] in_628,
  input [15:0] in_629,
  input [15:0] in_63,
  input [15:0] in_630,
  input [15:0] in_631,
  input [15:0] in_632,
  input [15:0] in_633,
  input [15:0] in_634,
  input [15:0] in_635,
  input [15:0] in_636,
  input [15:0] in_637,
  input [15:0] in_638,
  input [15:0] in_639,
  input [15:0] in_64,
  input [15:0] in_640,
  input [15:0] in_641,
  input [15:0] in_642,
  input [15:0] in_643,
  input [15:0] in_644,
  input [15:0] in_645,
  input [15:0] in_646,
  input [15:0] in_647,
  input [15:0] in_648,
  input [15:0] in_649,
  input [15:0] in_65,
  input [15:0] in_650,
  input [15:0] in_651,
  input [15:0] in_652,
  input [15:0] in_653,
  input [15:0] in_654,
  input [15:0] in_655,
  input [15:0] in_656,
  input [15:0] in_657,
  input [15:0] in_658,
  input [15:0] in_659,
  input [15:0] in_66,
  input [15:0] in_660,
  input [15:0] in_661,
  input [15:0] in_662,
  input [15:0] in_663,
  input [15:0] in_664,
  input [15:0] in_665,
  input [15:0] in_666,
  input [15:0] in_667,
  input [15:0] in_668,
  input [15:0] in_669,
  input [15:0] in_67,
  input [15:0] in_670,
  input [15:0] in_671,
  input [15:0] in_672,
  input [15:0] in_673,
  input [15:0] in_674,
  input [15:0] in_675,
  input [15:0] in_676,
  input [15:0] in_677,
  input [15:0] in_678,
  input [15:0] in_679,
  input [15:0] in_68,
  input [15:0] in_680,
  input [15:0] in_681,
  input [15:0] in_682,
  input [15:0] in_683,
  input [15:0] in_684,
  input [15:0] in_685,
  input [15:0] in_686,
  input [15:0] in_687,
  input [15:0] in_688,
  input [15:0] in_689,
  input [15:0] in_69,
  input [15:0] in_690,
  input [15:0] in_691,
  input [15:0] in_692,
  input [15:0] in_693,
  input [15:0] in_694,
  input [15:0] in_695,
  input [15:0] in_696,
  input [15:0] in_697,
  input [15:0] in_698,
  input [15:0] in_699,
  input [15:0] in_7,
  input [15:0] in_70,
  input [15:0] in_700,
  input [15:0] in_701,
  input [15:0] in_702,
  input [15:0] in_703,
  input [15:0] in_704,
  input [15:0] in_705,
  input [15:0] in_706,
  input [15:0] in_707,
  input [15:0] in_708,
  input [15:0] in_709,
  input [15:0] in_71,
  input [15:0] in_710,
  input [15:0] in_711,
  input [15:0] in_712,
  input [15:0] in_713,
  input [15:0] in_714,
  input [15:0] in_715,
  input [15:0] in_716,
  input [15:0] in_717,
  input [15:0] in_718,
  input [15:0] in_719,
  input [15:0] in_72,
  input [15:0] in_720,
  input [15:0] in_721,
  input [15:0] in_722,
  input [15:0] in_723,
  input [15:0] in_724,
  input [15:0] in_725,
  input [15:0] in_726,
  input [15:0] in_727,
  input [15:0] in_728,
  input [15:0] in_729,
  input [15:0] in_73,
  input [15:0] in_730,
  input [15:0] in_731,
  input [15:0] in_732,
  input [15:0] in_733,
  input [15:0] in_734,
  input [15:0] in_735,
  input [15:0] in_736,
  input [15:0] in_737,
  input [15:0] in_738,
  input [15:0] in_739,
  input [15:0] in_74,
  input [15:0] in_740,
  input [15:0] in_741,
  input [15:0] in_742,
  input [15:0] in_743,
  input [15:0] in_744,
  input [15:0] in_745,
  input [15:0] in_746,
  input [15:0] in_747,
  input [15:0] in_748,
  input [15:0] in_749,
  input [15:0] in_75,
  input [15:0] in_750,
  input [15:0] in_751,
  input [15:0] in_752,
  input [15:0] in_753,
  input [15:0] in_754,
  input [15:0] in_755,
  input [15:0] in_756,
  input [15:0] in_757,
  input [15:0] in_758,
  input [15:0] in_759,
  input [15:0] in_76,
  input [15:0] in_760,
  input [15:0] in_761,
  input [15:0] in_762,
  input [15:0] in_763,
  input [15:0] in_764,
  input [15:0] in_765,
  input [15:0] in_766,
  input [15:0] in_767,
  input [15:0] in_768,
  input [15:0] in_769,
  input [15:0] in_77,
  input [15:0] in_770,
  input [15:0] in_771,
  input [15:0] in_772,
  input [15:0] in_773,
  input [15:0] in_774,
  input [15:0] in_775,
  input [15:0] in_776,
  input [15:0] in_777,
  input [15:0] in_778,
  input [15:0] in_779,
  input [15:0] in_78,
  input [15:0] in_780,
  input [15:0] in_781,
  input [15:0] in_782,
  input [15:0] in_783,
  input [15:0] in_784,
  input [15:0] in_785,
  input [15:0] in_786,
  input [15:0] in_787,
  input [15:0] in_788,
  input [15:0] in_789,
  input [15:0] in_79,
  input [15:0] in_790,
  input [15:0] in_791,
  input [15:0] in_792,
  input [15:0] in_793,
  input [15:0] in_794,
  input [15:0] in_795,
  input [15:0] in_796,
  input [15:0] in_797,
  input [15:0] in_798,
  input [15:0] in_799,
  input [15:0] in_8,
  input [15:0] in_80,
  input [15:0] in_800,
  input [15:0] in_801,
  input [15:0] in_802,
  input [15:0] in_803,
  input [15:0] in_804,
  input [15:0] in_805,
  input [15:0] in_806,
  input [15:0] in_807,
  input [15:0] in_808,
  input [15:0] in_809,
  input [15:0] in_81,
  input [15:0] in_810,
  input [15:0] in_811,
  input [15:0] in_812,
  input [15:0] in_813,
  input [15:0] in_814,
  input [15:0] in_815,
  input [15:0] in_816,
  input [15:0] in_817,
  input [15:0] in_818,
  input [15:0] in_819,
  input [15:0] in_82,
  input [15:0] in_820,
  input [15:0] in_821,
  input [15:0] in_822,
  input [15:0] in_823,
  input [15:0] in_824,
  input [15:0] in_825,
  input [15:0] in_826,
  input [15:0] in_827,
  input [15:0] in_828,
  input [15:0] in_829,
  input [15:0] in_83,
  input [15:0] in_830,
  input [15:0] in_831,
  input [15:0] in_832,
  input [15:0] in_833,
  input [15:0] in_834,
  input [15:0] in_835,
  input [15:0] in_836,
  input [15:0] in_837,
  input [15:0] in_838,
  input [15:0] in_839,
  input [15:0] in_84,
  input [15:0] in_840,
  input [15:0] in_841,
  input [15:0] in_842,
  input [15:0] in_843,
  input [15:0] in_844,
  input [15:0] in_845,
  input [15:0] in_846,
  input [15:0] in_847,
  input [15:0] in_848,
  input [15:0] in_849,
  input [15:0] in_85,
  input [15:0] in_850,
  input [15:0] in_851,
  input [15:0] in_852,
  input [15:0] in_853,
  input [15:0] in_854,
  input [15:0] in_855,
  input [15:0] in_856,
  input [15:0] in_857,
  input [15:0] in_858,
  input [15:0] in_859,
  input [15:0] in_86,
  input [15:0] in_860,
  input [15:0] in_861,
  input [15:0] in_862,
  input [15:0] in_863,
  input [15:0] in_864,
  input [15:0] in_865,
  input [15:0] in_866,
  input [15:0] in_867,
  input [15:0] in_868,
  input [15:0] in_869,
  input [15:0] in_87,
  input [15:0] in_870,
  input [15:0] in_871,
  input [15:0] in_872,
  input [15:0] in_873,
  input [15:0] in_874,
  input [15:0] in_875,
  input [15:0] in_876,
  input [15:0] in_877,
  input [15:0] in_878,
  input [15:0] in_879,
  input [15:0] in_88,
  input [15:0] in_880,
  input [15:0] in_881,
  input [15:0] in_882,
  input [15:0] in_883,
  input [15:0] in_884,
  input [15:0] in_885,
  input [15:0] in_886,
  input [15:0] in_887,
  input [15:0] in_888,
  input [15:0] in_889,
  input [15:0] in_89,
  input [15:0] in_890,
  input [15:0] in_891,
  input [15:0] in_892,
  input [15:0] in_893,
  input [15:0] in_894,
  input [15:0] in_895,
  input [15:0] in_896,
  input [15:0] in_897,
  input [15:0] in_898,
  input [15:0] in_899,
  input [15:0] in_9,
  input [15:0] in_90,
  input [15:0] in_900,
  input [15:0] in_901,
  input [15:0] in_902,
  input [15:0] in_903,
  input [15:0] in_904,
  input [15:0] in_905,
  input [15:0] in_906,
  input [15:0] in_907,
  input [15:0] in_908,
  input [15:0] in_909,
  input [15:0] in_91,
  input [15:0] in_910,
  input [15:0] in_911,
  input [15:0] in_912,
  input [15:0] in_913,
  input [15:0] in_914,
  input [15:0] in_915,
  input [15:0] in_916,
  input [15:0] in_917,
  input [15:0] in_918,
  input [15:0] in_919,
  input [15:0] in_92,
  input [15:0] in_920,
  input [15:0] in_921,
  input [15:0] in_922,
  input [15:0] in_923,
  input [15:0] in_924,
  input [15:0] in_925,
  input [15:0] in_926,
  input [15:0] in_927,
  input [15:0] in_928,
  input [15:0] in_929,
  input [15:0] in_93,
  input [15:0] in_930,
  input [15:0] in_931,
  input [15:0] in_932,
  input [15:0] in_933,
  input [15:0] in_934,
  input [15:0] in_935,
  input [15:0] in_936,
  input [15:0] in_937,
  input [15:0] in_938,
  input [15:0] in_939,
  input [15:0] in_94,
  input [15:0] in_940,
  input [15:0] in_941,
  input [15:0] in_942,
  input [15:0] in_943,
  input [15:0] in_944,
  input [15:0] in_945,
  input [15:0] in_946,
  input [15:0] in_947,
  input [15:0] in_948,
  input [15:0] in_949,
  input [15:0] in_95,
  input [15:0] in_950,
  input [15:0] in_951,
  input [15:0] in_952,
  input [15:0] in_953,
  input [15:0] in_954,
  input [15:0] in_955,
  input [15:0] in_956,
  input [15:0] in_957,
  input [15:0] in_958,
  input [15:0] in_959,
  input [15:0] in_96,
  input [15:0] in_960,
  input [15:0] in_961,
  input [15:0] in_962,
  input [15:0] in_963,
  input [15:0] in_964,
  input [15:0] in_965,
  input [15:0] in_966,
  input [15:0] in_967,
  input [15:0] in_968,
  input [15:0] in_969,
  input [15:0] in_97,
  input [15:0] in_970,
  input [15:0] in_971,
  input [15:0] in_972,
  input [15:0] in_973,
  input [15:0] in_974,
  input [15:0] in_975,
  input [15:0] in_976,
  input [15:0] in_977,
  input [15:0] in_978,
  input [15:0] in_979,
  input [15:0] in_98,
  input [15:0] in_980,
  input [15:0] in_981,
  input [15:0] in_982,
  input [15:0] in_983,
  input [15:0] in_984,
  input [15:0] in_985,
  input [15:0] in_986,
  input [15:0] in_987,
  input [15:0] in_988,
  input [15:0] in_989,
  input [15:0] in_99,
  input [15:0] in_990,
  input [15:0] in_991,
  input [15:0] in_992,
  input [15:0] in_993,
  input [15:0] in_994,
  input [15:0] in_995,
  input [15:0] in_996,
  input [15:0] in_997,
  input [15:0] in_998,
  input [15:0] in_999,
  output [15:0] out_0,
  output [15:0] out_1,
  output [15:0] out_10,
  output [15:0] out_100,
  output [15:0] out_101,
  output [15:0] out_102,
  output [15:0] out_103,
  output [15:0] out_104,
  output [15:0] out_105,
  output [15:0] out_106,
  output [15:0] out_107,
  output [15:0] out_108,
  output [15:0] out_109,
  output [15:0] out_11,
  output [15:0] out_110,
  output [15:0] out_111,
  output [15:0] out_112,
  output [15:0] out_113,
  output [15:0] out_114,
  output [15:0] out_115,
  output [15:0] out_116,
  output [15:0] out_117,
  output [15:0] out_118,
  output [15:0] out_119,
  output [15:0] out_12,
  output [15:0] out_120,
  output [15:0] out_121,
  output [15:0] out_122,
  output [15:0] out_123,
  output [15:0] out_124,
  output [15:0] out_125,
  output [15:0] out_126,
  output [15:0] out_127,
  output [15:0] out_128,
  output [15:0] out_129,
  output [15:0] out_13,
  output [15:0] out_130,
  output [15:0] out_131,
  output [15:0] out_132,
  output [15:0] out_133,
  output [15:0] out_134,
  output [15:0] out_135,
  output [15:0] out_136,
  output [15:0] out_137,
  output [15:0] out_138,
  output [15:0] out_139,
  output [15:0] out_14,
  output [15:0] out_140,
  output [15:0] out_141,
  output [15:0] out_142,
  output [15:0] out_143,
  output [15:0] out_144,
  output [15:0] out_145,
  output [15:0] out_146,
  output [15:0] out_147,
  output [15:0] out_148,
  output [15:0] out_149,
  output [15:0] out_15,
  output [15:0] out_150,
  output [15:0] out_151,
  output [15:0] out_152,
  output [15:0] out_153,
  output [15:0] out_154,
  output [15:0] out_155,
  output [15:0] out_156,
  output [15:0] out_157,
  output [15:0] out_158,
  output [15:0] out_159,
  output [15:0] out_16,
  output [15:0] out_160,
  output [15:0] out_161,
  output [15:0] out_162,
  output [15:0] out_163,
  output [15:0] out_164,
  output [15:0] out_165,
  output [15:0] out_166,
  output [15:0] out_167,
  output [15:0] out_168,
  output [15:0] out_169,
  output [15:0] out_17,
  output [15:0] out_170,
  output [15:0] out_171,
  output [15:0] out_172,
  output [15:0] out_173,
  output [15:0] out_174,
  output [15:0] out_175,
  output [15:0] out_176,
  output [15:0] out_177,
  output [15:0] out_178,
  output [15:0] out_179,
  output [15:0] out_18,
  output [15:0] out_180,
  output [15:0] out_181,
  output [15:0] out_182,
  output [15:0] out_183,
  output [15:0] out_184,
  output [15:0] out_185,
  output [15:0] out_186,
  output [15:0] out_187,
  output [15:0] out_188,
  output [15:0] out_189,
  output [15:0] out_19,
  output [15:0] out_190,
  output [15:0] out_191,
  output [15:0] out_192,
  output [15:0] out_193,
  output [15:0] out_194,
  output [15:0] out_195,
  output [15:0] out_196,
  output [15:0] out_197,
  output [15:0] out_198,
  output [15:0] out_199,
  output [15:0] out_2,
  output [15:0] out_20,
  output [15:0] out_200,
  output [15:0] out_201,
  output [15:0] out_202,
  output [15:0] out_203,
  output [15:0] out_204,
  output [15:0] out_205,
  output [15:0] out_206,
  output [15:0] out_207,
  output [15:0] out_208,
  output [15:0] out_209,
  output [15:0] out_21,
  output [15:0] out_210,
  output [15:0] out_211,
  output [15:0] out_212,
  output [15:0] out_213,
  output [15:0] out_214,
  output [15:0] out_215,
  output [15:0] out_216,
  output [15:0] out_217,
  output [15:0] out_218,
  output [15:0] out_219,
  output [15:0] out_22,
  output [15:0] out_220,
  output [15:0] out_221,
  output [15:0] out_222,
  output [15:0] out_223,
  output [15:0] out_224,
  output [15:0] out_225,
  output [15:0] out_226,
  output [15:0] out_227,
  output [15:0] out_228,
  output [15:0] out_229,
  output [15:0] out_23,
  output [15:0] out_230,
  output [15:0] out_231,
  output [15:0] out_232,
  output [15:0] out_233,
  output [15:0] out_234,
  output [15:0] out_235,
  output [15:0] out_236,
  output [15:0] out_237,
  output [15:0] out_238,
  output [15:0] out_239,
  output [15:0] out_24,
  output [15:0] out_240,
  output [15:0] out_241,
  output [15:0] out_242,
  output [15:0] out_243,
  output [15:0] out_244,
  output [15:0] out_245,
  output [15:0] out_246,
  output [15:0] out_247,
  output [15:0] out_248,
  output [15:0] out_249,
  output [15:0] out_25,
  output [15:0] out_250,
  output [15:0] out_251,
  output [15:0] out_252,
  output [15:0] out_253,
  output [15:0] out_254,
  output [15:0] out_255,
  output [15:0] out_256,
  output [15:0] out_257,
  output [15:0] out_258,
  output [15:0] out_259,
  output [15:0] out_26,
  output [15:0] out_260,
  output [15:0] out_261,
  output [15:0] out_262,
  output [15:0] out_263,
  output [15:0] out_264,
  output [15:0] out_265,
  output [15:0] out_266,
  output [15:0] out_267,
  output [15:0] out_268,
  output [15:0] out_269,
  output [15:0] out_27,
  output [15:0] out_270,
  output [15:0] out_271,
  output [15:0] out_272,
  output [15:0] out_273,
  output [15:0] out_274,
  output [15:0] out_275,
  output [15:0] out_276,
  output [15:0] out_277,
  output [15:0] out_278,
  output [15:0] out_279,
  output [15:0] out_28,
  output [15:0] out_280,
  output [15:0] out_281,
  output [15:0] out_282,
  output [15:0] out_283,
  output [15:0] out_284,
  output [15:0] out_285,
  output [15:0] out_286,
  output [15:0] out_287,
  output [15:0] out_288,
  output [15:0] out_289,
  output [15:0] out_29,
  output [15:0] out_290,
  output [15:0] out_291,
  output [15:0] out_292,
  output [15:0] out_293,
  output [15:0] out_294,
  output [15:0] out_295,
  output [15:0] out_296,
  output [15:0] out_297,
  output [15:0] out_298,
  output [15:0] out_299,
  output [15:0] out_3,
  output [15:0] out_30,
  output [15:0] out_300,
  output [15:0] out_301,
  output [15:0] out_302,
  output [15:0] out_303,
  output [15:0] out_304,
  output [15:0] out_305,
  output [15:0] out_306,
  output [15:0] out_307,
  output [15:0] out_308,
  output [15:0] out_309,
  output [15:0] out_31,
  output [15:0] out_310,
  output [15:0] out_311,
  output [15:0] out_312,
  output [15:0] out_313,
  output [15:0] out_314,
  output [15:0] out_315,
  output [15:0] out_316,
  output [15:0] out_317,
  output [15:0] out_318,
  output [15:0] out_319,
  output [15:0] out_32,
  output [15:0] out_320,
  output [15:0] out_321,
  output [15:0] out_322,
  output [15:0] out_323,
  output [15:0] out_324,
  output [15:0] out_325,
  output [15:0] out_326,
  output [15:0] out_327,
  output [15:0] out_328,
  output [15:0] out_329,
  output [15:0] out_33,
  output [15:0] out_330,
  output [15:0] out_331,
  output [15:0] out_332,
  output [15:0] out_333,
  output [15:0] out_334,
  output [15:0] out_335,
  output [15:0] out_336,
  output [15:0] out_337,
  output [15:0] out_338,
  output [15:0] out_339,
  output [15:0] out_34,
  output [15:0] out_340,
  output [15:0] out_341,
  output [15:0] out_342,
  output [15:0] out_343,
  output [15:0] out_344,
  output [15:0] out_345,
  output [15:0] out_346,
  output [15:0] out_347,
  output [15:0] out_348,
  output [15:0] out_349,
  output [15:0] out_35,
  output [15:0] out_350,
  output [15:0] out_351,
  output [15:0] out_352,
  output [15:0] out_353,
  output [15:0] out_354,
  output [15:0] out_355,
  output [15:0] out_356,
  output [15:0] out_357,
  output [15:0] out_358,
  output [15:0] out_359,
  output [15:0] out_36,
  output [15:0] out_360,
  output [15:0] out_361,
  output [15:0] out_362,
  output [15:0] out_363,
  output [15:0] out_364,
  output [15:0] out_365,
  output [15:0] out_366,
  output [15:0] out_367,
  output [15:0] out_368,
  output [15:0] out_369,
  output [15:0] out_37,
  output [15:0] out_370,
  output [15:0] out_371,
  output [15:0] out_372,
  output [15:0] out_373,
  output [15:0] out_374,
  output [15:0] out_375,
  output [15:0] out_376,
  output [15:0] out_377,
  output [15:0] out_378,
  output [15:0] out_379,
  output [15:0] out_38,
  output [15:0] out_380,
  output [15:0] out_381,
  output [15:0] out_382,
  output [15:0] out_383,
  output [15:0] out_384,
  output [15:0] out_385,
  output [15:0] out_386,
  output [15:0] out_387,
  output [15:0] out_388,
  output [15:0] out_389,
  output [15:0] out_39,
  output [15:0] out_390,
  output [15:0] out_391,
  output [15:0] out_392,
  output [15:0] out_393,
  output [15:0] out_394,
  output [15:0] out_395,
  output [15:0] out_396,
  output [15:0] out_397,
  output [15:0] out_398,
  output [15:0] out_399,
  output [15:0] out_4,
  output [15:0] out_40,
  output [15:0] out_400,
  output [15:0] out_401,
  output [15:0] out_402,
  output [15:0] out_403,
  output [15:0] out_404,
  output [15:0] out_405,
  output [15:0] out_406,
  output [15:0] out_407,
  output [15:0] out_408,
  output [15:0] out_409,
  output [15:0] out_41,
  output [15:0] out_410,
  output [15:0] out_411,
  output [15:0] out_412,
  output [15:0] out_413,
  output [15:0] out_414,
  output [15:0] out_415,
  output [15:0] out_416,
  output [15:0] out_417,
  output [15:0] out_418,
  output [15:0] out_419,
  output [15:0] out_42,
  output [15:0] out_420,
  output [15:0] out_421,
  output [15:0] out_422,
  output [15:0] out_423,
  output [15:0] out_424,
  output [15:0] out_425,
  output [15:0] out_426,
  output [15:0] out_427,
  output [15:0] out_428,
  output [15:0] out_429,
  output [15:0] out_43,
  output [15:0] out_430,
  output [15:0] out_431,
  output [15:0] out_432,
  output [15:0] out_433,
  output [15:0] out_434,
  output [15:0] out_435,
  output [15:0] out_436,
  output [15:0] out_437,
  output [15:0] out_438,
  output [15:0] out_439,
  output [15:0] out_44,
  output [15:0] out_440,
  output [15:0] out_441,
  output [15:0] out_442,
  output [15:0] out_443,
  output [15:0] out_444,
  output [15:0] out_445,
  output [15:0] out_446,
  output [15:0] out_447,
  output [15:0] out_448,
  output [15:0] out_449,
  output [15:0] out_45,
  output [15:0] out_450,
  output [15:0] out_451,
  output [15:0] out_452,
  output [15:0] out_453,
  output [15:0] out_454,
  output [15:0] out_455,
  output [15:0] out_456,
  output [15:0] out_457,
  output [15:0] out_458,
  output [15:0] out_459,
  output [15:0] out_46,
  output [15:0] out_460,
  output [15:0] out_461,
  output [15:0] out_462,
  output [15:0] out_463,
  output [15:0] out_464,
  output [15:0] out_465,
  output [15:0] out_466,
  output [15:0] out_467,
  output [15:0] out_468,
  output [15:0] out_469,
  output [15:0] out_47,
  output [15:0] out_470,
  output [15:0] out_471,
  output [15:0] out_472,
  output [15:0] out_473,
  output [15:0] out_474,
  output [15:0] out_475,
  output [15:0] out_476,
  output [15:0] out_477,
  output [15:0] out_478,
  output [15:0] out_479,
  output [15:0] out_48,
  output [15:0] out_480,
  output [15:0] out_481,
  output [15:0] out_482,
  output [15:0] out_483,
  output [15:0] out_484,
  output [15:0] out_485,
  output [15:0] out_486,
  output [15:0] out_487,
  output [15:0] out_488,
  output [15:0] out_489,
  output [15:0] out_49,
  output [15:0] out_490,
  output [15:0] out_491,
  output [15:0] out_492,
  output [15:0] out_493,
  output [15:0] out_494,
  output [15:0] out_495,
  output [15:0] out_496,
  output [15:0] out_497,
  output [15:0] out_498,
  output [15:0] out_499,
  output [15:0] out_5,
  output [15:0] out_50,
  output [15:0] out_500,
  output [15:0] out_501,
  output [15:0] out_502,
  output [15:0] out_503,
  output [15:0] out_504,
  output [15:0] out_505,
  output [15:0] out_506,
  output [15:0] out_507,
  output [15:0] out_508,
  output [15:0] out_509,
  output [15:0] out_51,
  output [15:0] out_510,
  output [15:0] out_511,
  output [15:0] out_512,
  output [15:0] out_513,
  output [15:0] out_514,
  output [15:0] out_515,
  output [15:0] out_516,
  output [15:0] out_517,
  output [15:0] out_518,
  output [15:0] out_519,
  output [15:0] out_52,
  output [15:0] out_520,
  output [15:0] out_521,
  output [15:0] out_522,
  output [15:0] out_523,
  output [15:0] out_524,
  output [15:0] out_525,
  output [15:0] out_526,
  output [15:0] out_527,
  output [15:0] out_528,
  output [15:0] out_529,
  output [15:0] out_53,
  output [15:0] out_530,
  output [15:0] out_531,
  output [15:0] out_532,
  output [15:0] out_533,
  output [15:0] out_534,
  output [15:0] out_535,
  output [15:0] out_536,
  output [15:0] out_537,
  output [15:0] out_538,
  output [15:0] out_539,
  output [15:0] out_54,
  output [15:0] out_540,
  output [15:0] out_541,
  output [15:0] out_542,
  output [15:0] out_543,
  output [15:0] out_544,
  output [15:0] out_545,
  output [15:0] out_546,
  output [15:0] out_547,
  output [15:0] out_548,
  output [15:0] out_549,
  output [15:0] out_55,
  output [15:0] out_550,
  output [15:0] out_551,
  output [15:0] out_552,
  output [15:0] out_553,
  output [15:0] out_554,
  output [15:0] out_555,
  output [15:0] out_556,
  output [15:0] out_557,
  output [15:0] out_558,
  output [15:0] out_559,
  output [15:0] out_56,
  output [15:0] out_560,
  output [15:0] out_561,
  output [15:0] out_562,
  output [15:0] out_563,
  output [15:0] out_564,
  output [15:0] out_565,
  output [15:0] out_566,
  output [15:0] out_567,
  output [15:0] out_568,
  output [15:0] out_569,
  output [15:0] out_57,
  output [15:0] out_570,
  output [15:0] out_571,
  output [15:0] out_572,
  output [15:0] out_573,
  output [15:0] out_574,
  output [15:0] out_575,
  output [15:0] out_576,
  output [15:0] out_577,
  output [15:0] out_578,
  output [15:0] out_579,
  output [15:0] out_58,
  output [15:0] out_580,
  output [15:0] out_581,
  output [15:0] out_582,
  output [15:0] out_583,
  output [15:0] out_584,
  output [15:0] out_585,
  output [15:0] out_586,
  output [15:0] out_587,
  output [15:0] out_588,
  output [15:0] out_589,
  output [15:0] out_59,
  output [15:0] out_590,
  output [15:0] out_591,
  output [15:0] out_592,
  output [15:0] out_593,
  output [15:0] out_594,
  output [15:0] out_595,
  output [15:0] out_596,
  output [15:0] out_597,
  output [15:0] out_598,
  output [15:0] out_599,
  output [15:0] out_6,
  output [15:0] out_60,
  output [15:0] out_600,
  output [15:0] out_601,
  output [15:0] out_602,
  output [15:0] out_603,
  output [15:0] out_604,
  output [15:0] out_605,
  output [15:0] out_606,
  output [15:0] out_607,
  output [15:0] out_608,
  output [15:0] out_609,
  output [15:0] out_61,
  output [15:0] out_610,
  output [15:0] out_611,
  output [15:0] out_612,
  output [15:0] out_613,
  output [15:0] out_614,
  output [15:0] out_615,
  output [15:0] out_616,
  output [15:0] out_617,
  output [15:0] out_618,
  output [15:0] out_619,
  output [15:0] out_62,
  output [15:0] out_620,
  output [15:0] out_621,
  output [15:0] out_622,
  output [15:0] out_623,
  output [15:0] out_624,
  output [15:0] out_625,
  output [15:0] out_626,
  output [15:0] out_627,
  output [15:0] out_628,
  output [15:0] out_629,
  output [15:0] out_63,
  output [15:0] out_630,
  output [15:0] out_631,
  output [15:0] out_632,
  output [15:0] out_633,
  output [15:0] out_634,
  output [15:0] out_635,
  output [15:0] out_636,
  output [15:0] out_637,
  output [15:0] out_638,
  output [15:0] out_639,
  output [15:0] out_64,
  output [15:0] out_640,
  output [15:0] out_641,
  output [15:0] out_642,
  output [15:0] out_643,
  output [15:0] out_644,
  output [15:0] out_645,
  output [15:0] out_646,
  output [15:0] out_647,
  output [15:0] out_648,
  output [15:0] out_649,
  output [15:0] out_65,
  output [15:0] out_650,
  output [15:0] out_651,
  output [15:0] out_652,
  output [15:0] out_653,
  output [15:0] out_654,
  output [15:0] out_655,
  output [15:0] out_656,
  output [15:0] out_657,
  output [15:0] out_658,
  output [15:0] out_659,
  output [15:0] out_66,
  output [15:0] out_660,
  output [15:0] out_661,
  output [15:0] out_662,
  output [15:0] out_663,
  output [15:0] out_664,
  output [15:0] out_665,
  output [15:0] out_666,
  output [15:0] out_667,
  output [15:0] out_668,
  output [15:0] out_669,
  output [15:0] out_67,
  output [15:0] out_670,
  output [15:0] out_671,
  output [15:0] out_672,
  output [15:0] out_673,
  output [15:0] out_674,
  output [15:0] out_675,
  output [15:0] out_676,
  output [15:0] out_677,
  output [15:0] out_678,
  output [15:0] out_679,
  output [15:0] out_68,
  output [15:0] out_680,
  output [15:0] out_681,
  output [15:0] out_682,
  output [15:0] out_683,
  output [15:0] out_684,
  output [15:0] out_685,
  output [15:0] out_686,
  output [15:0] out_687,
  output [15:0] out_688,
  output [15:0] out_689,
  output [15:0] out_69,
  output [15:0] out_690,
  output [15:0] out_691,
  output [15:0] out_692,
  output [15:0] out_693,
  output [15:0] out_694,
  output [15:0] out_695,
  output [15:0] out_696,
  output [15:0] out_697,
  output [15:0] out_698,
  output [15:0] out_699,
  output [15:0] out_7,
  output [15:0] out_70,
  output [15:0] out_700,
  output [15:0] out_701,
  output [15:0] out_702,
  output [15:0] out_703,
  output [15:0] out_704,
  output [15:0] out_705,
  output [15:0] out_706,
  output [15:0] out_707,
  output [15:0] out_708,
  output [15:0] out_709,
  output [15:0] out_71,
  output [15:0] out_710,
  output [15:0] out_711,
  output [15:0] out_712,
  output [15:0] out_713,
  output [15:0] out_714,
  output [15:0] out_715,
  output [15:0] out_716,
  output [15:0] out_717,
  output [15:0] out_718,
  output [15:0] out_719,
  output [15:0] out_72,
  output [15:0] out_720,
  output [15:0] out_721,
  output [15:0] out_722,
  output [15:0] out_723,
  output [15:0] out_724,
  output [15:0] out_725,
  output [15:0] out_726,
  output [15:0] out_727,
  output [15:0] out_728,
  output [15:0] out_729,
  output [15:0] out_73,
  output [15:0] out_730,
  output [15:0] out_731,
  output [15:0] out_732,
  output [15:0] out_733,
  output [15:0] out_734,
  output [15:0] out_735,
  output [15:0] out_736,
  output [15:0] out_737,
  output [15:0] out_738,
  output [15:0] out_739,
  output [15:0] out_74,
  output [15:0] out_740,
  output [15:0] out_741,
  output [15:0] out_742,
  output [15:0] out_743,
  output [15:0] out_744,
  output [15:0] out_745,
  output [15:0] out_746,
  output [15:0] out_747,
  output [15:0] out_748,
  output [15:0] out_749,
  output [15:0] out_75,
  output [15:0] out_750,
  output [15:0] out_751,
  output [15:0] out_752,
  output [15:0] out_753,
  output [15:0] out_754,
  output [15:0] out_755,
  output [15:0] out_756,
  output [15:0] out_757,
  output [15:0] out_758,
  output [15:0] out_759,
  output [15:0] out_76,
  output [15:0] out_760,
  output [15:0] out_761,
  output [15:0] out_762,
  output [15:0] out_763,
  output [15:0] out_764,
  output [15:0] out_765,
  output [15:0] out_766,
  output [15:0] out_767,
  output [15:0] out_768,
  output [15:0] out_769,
  output [15:0] out_77,
  output [15:0] out_770,
  output [15:0] out_771,
  output [15:0] out_772,
  output [15:0] out_773,
  output [15:0] out_774,
  output [15:0] out_775,
  output [15:0] out_776,
  output [15:0] out_777,
  output [15:0] out_778,
  output [15:0] out_779,
  output [15:0] out_78,
  output [15:0] out_780,
  output [15:0] out_781,
  output [15:0] out_782,
  output [15:0] out_783,
  output [15:0] out_784,
  output [15:0] out_785,
  output [15:0] out_786,
  output [15:0] out_787,
  output [15:0] out_788,
  output [15:0] out_789,
  output [15:0] out_79,
  output [15:0] out_790,
  output [15:0] out_791,
  output [15:0] out_792,
  output [15:0] out_793,
  output [15:0] out_794,
  output [15:0] out_795,
  output [15:0] out_796,
  output [15:0] out_797,
  output [15:0] out_798,
  output [15:0] out_799,
  output [15:0] out_8,
  output [15:0] out_80,
  output [15:0] out_800,
  output [15:0] out_801,
  output [15:0] out_802,
  output [15:0] out_803,
  output [15:0] out_804,
  output [15:0] out_805,
  output [15:0] out_806,
  output [15:0] out_807,
  output [15:0] out_808,
  output [15:0] out_809,
  output [15:0] out_81,
  output [15:0] out_810,
  output [15:0] out_811,
  output [15:0] out_812,
  output [15:0] out_813,
  output [15:0] out_814,
  output [15:0] out_815,
  output [15:0] out_816,
  output [15:0] out_817,
  output [15:0] out_818,
  output [15:0] out_819,
  output [15:0] out_82,
  output [15:0] out_820,
  output [15:0] out_821,
  output [15:0] out_822,
  output [15:0] out_823,
  output [15:0] out_824,
  output [15:0] out_825,
  output [15:0] out_826,
  output [15:0] out_827,
  output [15:0] out_828,
  output [15:0] out_829,
  output [15:0] out_83,
  output [15:0] out_830,
  output [15:0] out_831,
  output [15:0] out_832,
  output [15:0] out_833,
  output [15:0] out_834,
  output [15:0] out_835,
  output [15:0] out_836,
  output [15:0] out_837,
  output [15:0] out_838,
  output [15:0] out_839,
  output [15:0] out_84,
  output [15:0] out_840,
  output [15:0] out_841,
  output [15:0] out_842,
  output [15:0] out_843,
  output [15:0] out_844,
  output [15:0] out_845,
  output [15:0] out_846,
  output [15:0] out_847,
  output [15:0] out_848,
  output [15:0] out_849,
  output [15:0] out_85,
  output [15:0] out_850,
  output [15:0] out_851,
  output [15:0] out_852,
  output [15:0] out_853,
  output [15:0] out_854,
  output [15:0] out_855,
  output [15:0] out_856,
  output [15:0] out_857,
  output [15:0] out_858,
  output [15:0] out_859,
  output [15:0] out_86,
  output [15:0] out_860,
  output [15:0] out_861,
  output [15:0] out_862,
  output [15:0] out_863,
  output [15:0] out_864,
  output [15:0] out_865,
  output [15:0] out_866,
  output [15:0] out_867,
  output [15:0] out_868,
  output [15:0] out_869,
  output [15:0] out_87,
  output [15:0] out_870,
  output [15:0] out_871,
  output [15:0] out_872,
  output [15:0] out_873,
  output [15:0] out_874,
  output [15:0] out_875,
  output [15:0] out_876,
  output [15:0] out_877,
  output [15:0] out_878,
  output [15:0] out_879,
  output [15:0] out_88,
  output [15:0] out_880,
  output [15:0] out_881,
  output [15:0] out_882,
  output [15:0] out_883,
  output [15:0] out_884,
  output [15:0] out_885,
  output [15:0] out_886,
  output [15:0] out_887,
  output [15:0] out_888,
  output [15:0] out_889,
  output [15:0] out_89,
  output [15:0] out_890,
  output [15:0] out_891,
  output [15:0] out_892,
  output [15:0] out_893,
  output [15:0] out_894,
  output [15:0] out_895,
  output [15:0] out_896,
  output [15:0] out_897,
  output [15:0] out_898,
  output [15:0] out_899,
  output [15:0] out_9,
  output [15:0] out_90,
  output [15:0] out_900,
  output [15:0] out_901,
  output [15:0] out_902,
  output [15:0] out_903,
  output [15:0] out_904,
  output [15:0] out_905,
  output [15:0] out_906,
  output [15:0] out_907,
  output [15:0] out_908,
  output [15:0] out_909,
  output [15:0] out_91,
  output [15:0] out_910,
  output [15:0] out_911,
  output [15:0] out_912,
  output [15:0] out_913,
  output [15:0] out_914,
  output [15:0] out_915,
  output [15:0] out_916,
  output [15:0] out_917,
  output [15:0] out_918,
  output [15:0] out_919,
  output [15:0] out_92,
  output [15:0] out_920,
  output [15:0] out_921,
  output [15:0] out_922,
  output [15:0] out_923,
  output [15:0] out_924,
  output [15:0] out_925,
  output [15:0] out_926,
  output [15:0] out_927,
  output [15:0] out_928,
  output [15:0] out_929,
  output [15:0] out_93,
  output [15:0] out_930,
  output [15:0] out_931,
  output [15:0] out_932,
  output [15:0] out_933,
  output [15:0] out_934,
  output [15:0] out_935,
  output [15:0] out_936,
  output [15:0] out_937,
  output [15:0] out_938,
  output [15:0] out_939,
  output [15:0] out_94,
  output [15:0] out_940,
  output [15:0] out_941,
  output [15:0] out_942,
  output [15:0] out_943,
  output [15:0] out_944,
  output [15:0] out_945,
  output [15:0] out_946,
  output [15:0] out_947,
  output [15:0] out_948,
  output [15:0] out_949,
  output [15:0] out_95,
  output [15:0] out_950,
  output [15:0] out_951,
  output [15:0] out_952,
  output [15:0] out_953,
  output [15:0] out_954,
  output [15:0] out_955,
  output [15:0] out_956,
  output [15:0] out_957,
  output [15:0] out_958,
  output [15:0] out_959,
  output [15:0] out_96,
  output [15:0] out_960,
  output [15:0] out_961,
  output [15:0] out_962,
  output [15:0] out_963,
  output [15:0] out_964,
  output [15:0] out_965,
  output [15:0] out_966,
  output [15:0] out_967,
  output [15:0] out_968,
  output [15:0] out_969,
  output [15:0] out_97,
  output [15:0] out_970,
  output [15:0] out_971,
  output [15:0] out_972,
  output [15:0] out_973,
  output [15:0] out_974,
  output [15:0] out_975,
  output [15:0] out_976,
  output [15:0] out_977,
  output [15:0] out_978,
  output [15:0] out_979,
  output [15:0] out_98,
  output [15:0] out_980,
  output [15:0] out_981,
  output [15:0] out_982,
  output [15:0] out_983,
  output [15:0] out_984,
  output [15:0] out_985,
  output [15:0] out_986,
  output [15:0] out_987,
  output [15:0] out_988,
  output [15:0] out_989,
  output [15:0] out_99,
  output [15:0] out_990,
  output [15:0] out_991,
  output [15:0] out_992,
  output [15:0] out_993,
  output [15:0] out_994,
  output [15:0] out_995,
  output [15:0] out_996,
  output [15:0] out_997,
  output [15:0] out_998,
  output [15:0] out_999
);
  //Wire declarations for instance 'and_0' (Module coreir_and)
  wire [15:0] and_0__in0;
  wire [15:0] and_0__in1;
  wire [15:0] and_0__out;
  coreir_and #(.width(16)) and_0(
    .in0(and_0__in0),
    .in1(and_0__in1),
    .out(and_0__out)
  );

  //Wire declarations for instance 'and_10' (Module coreir_and)
  wire [15:0] and_10__in0;
  wire [15:0] and_10__in1;
  wire [15:0] and_10__out;
  coreir_and #(.width(16)) and_10(
    .in0(and_10__in0),
    .in1(and_10__in1),
    .out(and_10__out)
  );

  //Wire declarations for instance 'and_100' (Module coreir_and)
  wire [15:0] and_100__in0;
  wire [15:0] and_100__in1;
  wire [15:0] and_100__out;
  coreir_and #(.width(16)) and_100(
    .in0(and_100__in0),
    .in1(and_100__in1),
    .out(and_100__out)
  );

  //Wire declarations for instance 'and_102' (Module coreir_and)
  wire [15:0] and_102__in0;
  wire [15:0] and_102__in1;
  wire [15:0] and_102__out;
  coreir_and #(.width(16)) and_102(
    .in0(and_102__in0),
    .in1(and_102__in1),
    .out(and_102__out)
  );

  //Wire declarations for instance 'and_104' (Module coreir_and)
  wire [15:0] and_104__in0;
  wire [15:0] and_104__in1;
  wire [15:0] and_104__out;
  coreir_and #(.width(16)) and_104(
    .in0(and_104__in0),
    .in1(and_104__in1),
    .out(and_104__out)
  );

  //Wire declarations for instance 'and_106' (Module coreir_and)
  wire [15:0] and_106__in0;
  wire [15:0] and_106__in1;
  wire [15:0] and_106__out;
  coreir_and #(.width(16)) and_106(
    .in0(and_106__in0),
    .in1(and_106__in1),
    .out(and_106__out)
  );

  //Wire declarations for instance 'and_108' (Module coreir_and)
  wire [15:0] and_108__in0;
  wire [15:0] and_108__in1;
  wire [15:0] and_108__out;
  coreir_and #(.width(16)) and_108(
    .in0(and_108__in0),
    .in1(and_108__in1),
    .out(and_108__out)
  );

  //Wire declarations for instance 'and_110' (Module coreir_and)
  wire [15:0] and_110__in0;
  wire [15:0] and_110__in1;
  wire [15:0] and_110__out;
  coreir_and #(.width(16)) and_110(
    .in0(and_110__in0),
    .in1(and_110__in1),
    .out(and_110__out)
  );

  //Wire declarations for instance 'and_112' (Module coreir_and)
  wire [15:0] and_112__in0;
  wire [15:0] and_112__in1;
  wire [15:0] and_112__out;
  coreir_and #(.width(16)) and_112(
    .in0(and_112__in0),
    .in1(and_112__in1),
    .out(and_112__out)
  );

  //Wire declarations for instance 'and_114' (Module coreir_and)
  wire [15:0] and_114__in0;
  wire [15:0] and_114__in1;
  wire [15:0] and_114__out;
  coreir_and #(.width(16)) and_114(
    .in0(and_114__in0),
    .in1(and_114__in1),
    .out(and_114__out)
  );

  //Wire declarations for instance 'and_116' (Module coreir_and)
  wire [15:0] and_116__in0;
  wire [15:0] and_116__in1;
  wire [15:0] and_116__out;
  coreir_and #(.width(16)) and_116(
    .in0(and_116__in0),
    .in1(and_116__in1),
    .out(and_116__out)
  );

  //Wire declarations for instance 'and_118' (Module coreir_and)
  wire [15:0] and_118__in0;
  wire [15:0] and_118__in1;
  wire [15:0] and_118__out;
  coreir_and #(.width(16)) and_118(
    .in0(and_118__in0),
    .in1(and_118__in1),
    .out(and_118__out)
  );

  //Wire declarations for instance 'and_12' (Module coreir_and)
  wire [15:0] and_12__in0;
  wire [15:0] and_12__in1;
  wire [15:0] and_12__out;
  coreir_and #(.width(16)) and_12(
    .in0(and_12__in0),
    .in1(and_12__in1),
    .out(and_12__out)
  );

  //Wire declarations for instance 'and_120' (Module coreir_and)
  wire [15:0] and_120__in0;
  wire [15:0] and_120__in1;
  wire [15:0] and_120__out;
  coreir_and #(.width(16)) and_120(
    .in0(and_120__in0),
    .in1(and_120__in1),
    .out(and_120__out)
  );

  //Wire declarations for instance 'and_122' (Module coreir_and)
  wire [15:0] and_122__in0;
  wire [15:0] and_122__in1;
  wire [15:0] and_122__out;
  coreir_and #(.width(16)) and_122(
    .in0(and_122__in0),
    .in1(and_122__in1),
    .out(and_122__out)
  );

  //Wire declarations for instance 'and_124' (Module coreir_and)
  wire [15:0] and_124__in0;
  wire [15:0] and_124__in1;
  wire [15:0] and_124__out;
  coreir_and #(.width(16)) and_124(
    .in0(and_124__in0),
    .in1(and_124__in1),
    .out(and_124__out)
  );

  //Wire declarations for instance 'and_126' (Module coreir_and)
  wire [15:0] and_126__in0;
  wire [15:0] and_126__in1;
  wire [15:0] and_126__out;
  coreir_and #(.width(16)) and_126(
    .in0(and_126__in0),
    .in1(and_126__in1),
    .out(and_126__out)
  );

  //Wire declarations for instance 'and_128' (Module coreir_and)
  wire [15:0] and_128__in0;
  wire [15:0] and_128__in1;
  wire [15:0] and_128__out;
  coreir_and #(.width(16)) and_128(
    .in0(and_128__in0),
    .in1(and_128__in1),
    .out(and_128__out)
  );

  //Wire declarations for instance 'and_130' (Module coreir_and)
  wire [15:0] and_130__in0;
  wire [15:0] and_130__in1;
  wire [15:0] and_130__out;
  coreir_and #(.width(16)) and_130(
    .in0(and_130__in0),
    .in1(and_130__in1),
    .out(and_130__out)
  );

  //Wire declarations for instance 'and_132' (Module coreir_and)
  wire [15:0] and_132__in0;
  wire [15:0] and_132__in1;
  wire [15:0] and_132__out;
  coreir_and #(.width(16)) and_132(
    .in0(and_132__in0),
    .in1(and_132__in1),
    .out(and_132__out)
  );

  //Wire declarations for instance 'and_134' (Module coreir_and)
  wire [15:0] and_134__in0;
  wire [15:0] and_134__in1;
  wire [15:0] and_134__out;
  coreir_and #(.width(16)) and_134(
    .in0(and_134__in0),
    .in1(and_134__in1),
    .out(and_134__out)
  );

  //Wire declarations for instance 'and_136' (Module coreir_and)
  wire [15:0] and_136__in0;
  wire [15:0] and_136__in1;
  wire [15:0] and_136__out;
  coreir_and #(.width(16)) and_136(
    .in0(and_136__in0),
    .in1(and_136__in1),
    .out(and_136__out)
  );

  //Wire declarations for instance 'and_138' (Module coreir_and)
  wire [15:0] and_138__in0;
  wire [15:0] and_138__in1;
  wire [15:0] and_138__out;
  coreir_and #(.width(16)) and_138(
    .in0(and_138__in0),
    .in1(and_138__in1),
    .out(and_138__out)
  );

  //Wire declarations for instance 'and_14' (Module coreir_and)
  wire [15:0] and_14__in0;
  wire [15:0] and_14__in1;
  wire [15:0] and_14__out;
  coreir_and #(.width(16)) and_14(
    .in0(and_14__in0),
    .in1(and_14__in1),
    .out(and_14__out)
  );

  //Wire declarations for instance 'and_140' (Module coreir_and)
  wire [15:0] and_140__in0;
  wire [15:0] and_140__in1;
  wire [15:0] and_140__out;
  coreir_and #(.width(16)) and_140(
    .in0(and_140__in0),
    .in1(and_140__in1),
    .out(and_140__out)
  );

  //Wire declarations for instance 'and_142' (Module coreir_and)
  wire [15:0] and_142__in0;
  wire [15:0] and_142__in1;
  wire [15:0] and_142__out;
  coreir_and #(.width(16)) and_142(
    .in0(and_142__in0),
    .in1(and_142__in1),
    .out(and_142__out)
  );

  //Wire declarations for instance 'and_144' (Module coreir_and)
  wire [15:0] and_144__in0;
  wire [15:0] and_144__in1;
  wire [15:0] and_144__out;
  coreir_and #(.width(16)) and_144(
    .in0(and_144__in0),
    .in1(and_144__in1),
    .out(and_144__out)
  );

  //Wire declarations for instance 'and_146' (Module coreir_and)
  wire [15:0] and_146__in0;
  wire [15:0] and_146__in1;
  wire [15:0] and_146__out;
  coreir_and #(.width(16)) and_146(
    .in0(and_146__in0),
    .in1(and_146__in1),
    .out(and_146__out)
  );

  //Wire declarations for instance 'and_148' (Module coreir_and)
  wire [15:0] and_148__in0;
  wire [15:0] and_148__in1;
  wire [15:0] and_148__out;
  coreir_and #(.width(16)) and_148(
    .in0(and_148__in0),
    .in1(and_148__in1),
    .out(and_148__out)
  );

  //Wire declarations for instance 'and_150' (Module coreir_and)
  wire [15:0] and_150__in0;
  wire [15:0] and_150__in1;
  wire [15:0] and_150__out;
  coreir_and #(.width(16)) and_150(
    .in0(and_150__in0),
    .in1(and_150__in1),
    .out(and_150__out)
  );

  //Wire declarations for instance 'and_152' (Module coreir_and)
  wire [15:0] and_152__in0;
  wire [15:0] and_152__in1;
  wire [15:0] and_152__out;
  coreir_and #(.width(16)) and_152(
    .in0(and_152__in0),
    .in1(and_152__in1),
    .out(and_152__out)
  );

  //Wire declarations for instance 'and_154' (Module coreir_and)
  wire [15:0] and_154__in0;
  wire [15:0] and_154__in1;
  wire [15:0] and_154__out;
  coreir_and #(.width(16)) and_154(
    .in0(and_154__in0),
    .in1(and_154__in1),
    .out(and_154__out)
  );

  //Wire declarations for instance 'and_156' (Module coreir_and)
  wire [15:0] and_156__in0;
  wire [15:0] and_156__in1;
  wire [15:0] and_156__out;
  coreir_and #(.width(16)) and_156(
    .in0(and_156__in0),
    .in1(and_156__in1),
    .out(and_156__out)
  );

  //Wire declarations for instance 'and_158' (Module coreir_and)
  wire [15:0] and_158__in0;
  wire [15:0] and_158__in1;
  wire [15:0] and_158__out;
  coreir_and #(.width(16)) and_158(
    .in0(and_158__in0),
    .in1(and_158__in1),
    .out(and_158__out)
  );

  //Wire declarations for instance 'and_16' (Module coreir_and)
  wire [15:0] and_16__in0;
  wire [15:0] and_16__in1;
  wire [15:0] and_16__out;
  coreir_and #(.width(16)) and_16(
    .in0(and_16__in0),
    .in1(and_16__in1),
    .out(and_16__out)
  );

  //Wire declarations for instance 'and_160' (Module coreir_and)
  wire [15:0] and_160__in0;
  wire [15:0] and_160__in1;
  wire [15:0] and_160__out;
  coreir_and #(.width(16)) and_160(
    .in0(and_160__in0),
    .in1(and_160__in1),
    .out(and_160__out)
  );

  //Wire declarations for instance 'and_162' (Module coreir_and)
  wire [15:0] and_162__in0;
  wire [15:0] and_162__in1;
  wire [15:0] and_162__out;
  coreir_and #(.width(16)) and_162(
    .in0(and_162__in0),
    .in1(and_162__in1),
    .out(and_162__out)
  );

  //Wire declarations for instance 'and_164' (Module coreir_and)
  wire [15:0] and_164__in0;
  wire [15:0] and_164__in1;
  wire [15:0] and_164__out;
  coreir_and #(.width(16)) and_164(
    .in0(and_164__in0),
    .in1(and_164__in1),
    .out(and_164__out)
  );

  //Wire declarations for instance 'and_166' (Module coreir_and)
  wire [15:0] and_166__in0;
  wire [15:0] and_166__in1;
  wire [15:0] and_166__out;
  coreir_and #(.width(16)) and_166(
    .in0(and_166__in0),
    .in1(and_166__in1),
    .out(and_166__out)
  );

  //Wire declarations for instance 'and_168' (Module coreir_and)
  wire [15:0] and_168__in0;
  wire [15:0] and_168__in1;
  wire [15:0] and_168__out;
  coreir_and #(.width(16)) and_168(
    .in0(and_168__in0),
    .in1(and_168__in1),
    .out(and_168__out)
  );

  //Wire declarations for instance 'and_170' (Module coreir_and)
  wire [15:0] and_170__in0;
  wire [15:0] and_170__in1;
  wire [15:0] and_170__out;
  coreir_and #(.width(16)) and_170(
    .in0(and_170__in0),
    .in1(and_170__in1),
    .out(and_170__out)
  );

  //Wire declarations for instance 'and_172' (Module coreir_and)
  wire [15:0] and_172__in0;
  wire [15:0] and_172__in1;
  wire [15:0] and_172__out;
  coreir_and #(.width(16)) and_172(
    .in0(and_172__in0),
    .in1(and_172__in1),
    .out(and_172__out)
  );

  //Wire declarations for instance 'and_174' (Module coreir_and)
  wire [15:0] and_174__in0;
  wire [15:0] and_174__in1;
  wire [15:0] and_174__out;
  coreir_and #(.width(16)) and_174(
    .in0(and_174__in0),
    .in1(and_174__in1),
    .out(and_174__out)
  );

  //Wire declarations for instance 'and_176' (Module coreir_and)
  wire [15:0] and_176__in0;
  wire [15:0] and_176__in1;
  wire [15:0] and_176__out;
  coreir_and #(.width(16)) and_176(
    .in0(and_176__in0),
    .in1(and_176__in1),
    .out(and_176__out)
  );

  //Wire declarations for instance 'and_178' (Module coreir_and)
  wire [15:0] and_178__in0;
  wire [15:0] and_178__in1;
  wire [15:0] and_178__out;
  coreir_and #(.width(16)) and_178(
    .in0(and_178__in0),
    .in1(and_178__in1),
    .out(and_178__out)
  );

  //Wire declarations for instance 'and_18' (Module coreir_and)
  wire [15:0] and_18__in0;
  wire [15:0] and_18__in1;
  wire [15:0] and_18__out;
  coreir_and #(.width(16)) and_18(
    .in0(and_18__in0),
    .in1(and_18__in1),
    .out(and_18__out)
  );

  //Wire declarations for instance 'and_180' (Module coreir_and)
  wire [15:0] and_180__in0;
  wire [15:0] and_180__in1;
  wire [15:0] and_180__out;
  coreir_and #(.width(16)) and_180(
    .in0(and_180__in0),
    .in1(and_180__in1),
    .out(and_180__out)
  );

  //Wire declarations for instance 'and_182' (Module coreir_and)
  wire [15:0] and_182__in0;
  wire [15:0] and_182__in1;
  wire [15:0] and_182__out;
  coreir_and #(.width(16)) and_182(
    .in0(and_182__in0),
    .in1(and_182__in1),
    .out(and_182__out)
  );

  //Wire declarations for instance 'and_184' (Module coreir_and)
  wire [15:0] and_184__in0;
  wire [15:0] and_184__in1;
  wire [15:0] and_184__out;
  coreir_and #(.width(16)) and_184(
    .in0(and_184__in0),
    .in1(and_184__in1),
    .out(and_184__out)
  );

  //Wire declarations for instance 'and_186' (Module coreir_and)
  wire [15:0] and_186__in0;
  wire [15:0] and_186__in1;
  wire [15:0] and_186__out;
  coreir_and #(.width(16)) and_186(
    .in0(and_186__in0),
    .in1(and_186__in1),
    .out(and_186__out)
  );

  //Wire declarations for instance 'and_188' (Module coreir_and)
  wire [15:0] and_188__in0;
  wire [15:0] and_188__in1;
  wire [15:0] and_188__out;
  coreir_and #(.width(16)) and_188(
    .in0(and_188__in0),
    .in1(and_188__in1),
    .out(and_188__out)
  );

  //Wire declarations for instance 'and_190' (Module coreir_and)
  wire [15:0] and_190__in0;
  wire [15:0] and_190__in1;
  wire [15:0] and_190__out;
  coreir_and #(.width(16)) and_190(
    .in0(and_190__in0),
    .in1(and_190__in1),
    .out(and_190__out)
  );

  //Wire declarations for instance 'and_192' (Module coreir_and)
  wire [15:0] and_192__in0;
  wire [15:0] and_192__in1;
  wire [15:0] and_192__out;
  coreir_and #(.width(16)) and_192(
    .in0(and_192__in0),
    .in1(and_192__in1),
    .out(and_192__out)
  );

  //Wire declarations for instance 'and_194' (Module coreir_and)
  wire [15:0] and_194__in0;
  wire [15:0] and_194__in1;
  wire [15:0] and_194__out;
  coreir_and #(.width(16)) and_194(
    .in0(and_194__in0),
    .in1(and_194__in1),
    .out(and_194__out)
  );

  //Wire declarations for instance 'and_196' (Module coreir_and)
  wire [15:0] and_196__in0;
  wire [15:0] and_196__in1;
  wire [15:0] and_196__out;
  coreir_and #(.width(16)) and_196(
    .in0(and_196__in0),
    .in1(and_196__in1),
    .out(and_196__out)
  );

  //Wire declarations for instance 'and_198' (Module coreir_and)
  wire [15:0] and_198__in0;
  wire [15:0] and_198__in1;
  wire [15:0] and_198__out;
  coreir_and #(.width(16)) and_198(
    .in0(and_198__in0),
    .in1(and_198__in1),
    .out(and_198__out)
  );

  //Wire declarations for instance 'and_2' (Module coreir_and)
  wire [15:0] and_2__in0;
  wire [15:0] and_2__in1;
  wire [15:0] and_2__out;
  coreir_and #(.width(16)) and_2(
    .in0(and_2__in0),
    .in1(and_2__in1),
    .out(and_2__out)
  );

  //Wire declarations for instance 'and_20' (Module coreir_and)
  wire [15:0] and_20__in0;
  wire [15:0] and_20__in1;
  wire [15:0] and_20__out;
  coreir_and #(.width(16)) and_20(
    .in0(and_20__in0),
    .in1(and_20__in1),
    .out(and_20__out)
  );

  //Wire declarations for instance 'and_200' (Module coreir_and)
  wire [15:0] and_200__in0;
  wire [15:0] and_200__in1;
  wire [15:0] and_200__out;
  coreir_and #(.width(16)) and_200(
    .in0(and_200__in0),
    .in1(and_200__in1),
    .out(and_200__out)
  );

  //Wire declarations for instance 'and_202' (Module coreir_and)
  wire [15:0] and_202__in0;
  wire [15:0] and_202__in1;
  wire [15:0] and_202__out;
  coreir_and #(.width(16)) and_202(
    .in0(and_202__in0),
    .in1(and_202__in1),
    .out(and_202__out)
  );

  //Wire declarations for instance 'and_204' (Module coreir_and)
  wire [15:0] and_204__in0;
  wire [15:0] and_204__in1;
  wire [15:0] and_204__out;
  coreir_and #(.width(16)) and_204(
    .in0(and_204__in0),
    .in1(and_204__in1),
    .out(and_204__out)
  );

  //Wire declarations for instance 'and_206' (Module coreir_and)
  wire [15:0] and_206__in0;
  wire [15:0] and_206__in1;
  wire [15:0] and_206__out;
  coreir_and #(.width(16)) and_206(
    .in0(and_206__in0),
    .in1(and_206__in1),
    .out(and_206__out)
  );

  //Wire declarations for instance 'and_208' (Module coreir_and)
  wire [15:0] and_208__in0;
  wire [15:0] and_208__in1;
  wire [15:0] and_208__out;
  coreir_and #(.width(16)) and_208(
    .in0(and_208__in0),
    .in1(and_208__in1),
    .out(and_208__out)
  );

  //Wire declarations for instance 'and_210' (Module coreir_and)
  wire [15:0] and_210__in0;
  wire [15:0] and_210__in1;
  wire [15:0] and_210__out;
  coreir_and #(.width(16)) and_210(
    .in0(and_210__in0),
    .in1(and_210__in1),
    .out(and_210__out)
  );

  //Wire declarations for instance 'and_212' (Module coreir_and)
  wire [15:0] and_212__in0;
  wire [15:0] and_212__in1;
  wire [15:0] and_212__out;
  coreir_and #(.width(16)) and_212(
    .in0(and_212__in0),
    .in1(and_212__in1),
    .out(and_212__out)
  );

  //Wire declarations for instance 'and_214' (Module coreir_and)
  wire [15:0] and_214__in0;
  wire [15:0] and_214__in1;
  wire [15:0] and_214__out;
  coreir_and #(.width(16)) and_214(
    .in0(and_214__in0),
    .in1(and_214__in1),
    .out(and_214__out)
  );

  //Wire declarations for instance 'and_216' (Module coreir_and)
  wire [15:0] and_216__in0;
  wire [15:0] and_216__in1;
  wire [15:0] and_216__out;
  coreir_and #(.width(16)) and_216(
    .in0(and_216__in0),
    .in1(and_216__in1),
    .out(and_216__out)
  );

  //Wire declarations for instance 'and_218' (Module coreir_and)
  wire [15:0] and_218__in0;
  wire [15:0] and_218__in1;
  wire [15:0] and_218__out;
  coreir_and #(.width(16)) and_218(
    .in0(and_218__in0),
    .in1(and_218__in1),
    .out(and_218__out)
  );

  //Wire declarations for instance 'and_22' (Module coreir_and)
  wire [15:0] and_22__in0;
  wire [15:0] and_22__in1;
  wire [15:0] and_22__out;
  coreir_and #(.width(16)) and_22(
    .in0(and_22__in0),
    .in1(and_22__in1),
    .out(and_22__out)
  );

  //Wire declarations for instance 'and_220' (Module coreir_and)
  wire [15:0] and_220__in0;
  wire [15:0] and_220__in1;
  wire [15:0] and_220__out;
  coreir_and #(.width(16)) and_220(
    .in0(and_220__in0),
    .in1(and_220__in1),
    .out(and_220__out)
  );

  //Wire declarations for instance 'and_222' (Module coreir_and)
  wire [15:0] and_222__in0;
  wire [15:0] and_222__in1;
  wire [15:0] and_222__out;
  coreir_and #(.width(16)) and_222(
    .in0(and_222__in0),
    .in1(and_222__in1),
    .out(and_222__out)
  );

  //Wire declarations for instance 'and_224' (Module coreir_and)
  wire [15:0] and_224__in0;
  wire [15:0] and_224__in1;
  wire [15:0] and_224__out;
  coreir_and #(.width(16)) and_224(
    .in0(and_224__in0),
    .in1(and_224__in1),
    .out(and_224__out)
  );

  //Wire declarations for instance 'and_226' (Module coreir_and)
  wire [15:0] and_226__in0;
  wire [15:0] and_226__in1;
  wire [15:0] and_226__out;
  coreir_and #(.width(16)) and_226(
    .in0(and_226__in0),
    .in1(and_226__in1),
    .out(and_226__out)
  );

  //Wire declarations for instance 'and_228' (Module coreir_and)
  wire [15:0] and_228__in0;
  wire [15:0] and_228__in1;
  wire [15:0] and_228__out;
  coreir_and #(.width(16)) and_228(
    .in0(and_228__in0),
    .in1(and_228__in1),
    .out(and_228__out)
  );

  //Wire declarations for instance 'and_230' (Module coreir_and)
  wire [15:0] and_230__in0;
  wire [15:0] and_230__in1;
  wire [15:0] and_230__out;
  coreir_and #(.width(16)) and_230(
    .in0(and_230__in0),
    .in1(and_230__in1),
    .out(and_230__out)
  );

  //Wire declarations for instance 'and_232' (Module coreir_and)
  wire [15:0] and_232__in0;
  wire [15:0] and_232__in1;
  wire [15:0] and_232__out;
  coreir_and #(.width(16)) and_232(
    .in0(and_232__in0),
    .in1(and_232__in1),
    .out(and_232__out)
  );

  //Wire declarations for instance 'and_234' (Module coreir_and)
  wire [15:0] and_234__in0;
  wire [15:0] and_234__in1;
  wire [15:0] and_234__out;
  coreir_and #(.width(16)) and_234(
    .in0(and_234__in0),
    .in1(and_234__in1),
    .out(and_234__out)
  );

  //Wire declarations for instance 'and_236' (Module coreir_and)
  wire [15:0] and_236__in0;
  wire [15:0] and_236__in1;
  wire [15:0] and_236__out;
  coreir_and #(.width(16)) and_236(
    .in0(and_236__in0),
    .in1(and_236__in1),
    .out(and_236__out)
  );

  //Wire declarations for instance 'and_238' (Module coreir_and)
  wire [15:0] and_238__in0;
  wire [15:0] and_238__in1;
  wire [15:0] and_238__out;
  coreir_and #(.width(16)) and_238(
    .in0(and_238__in0),
    .in1(and_238__in1),
    .out(and_238__out)
  );

  //Wire declarations for instance 'and_24' (Module coreir_and)
  wire [15:0] and_24__in0;
  wire [15:0] and_24__in1;
  wire [15:0] and_24__out;
  coreir_and #(.width(16)) and_24(
    .in0(and_24__in0),
    .in1(and_24__in1),
    .out(and_24__out)
  );

  //Wire declarations for instance 'and_240' (Module coreir_and)
  wire [15:0] and_240__in0;
  wire [15:0] and_240__in1;
  wire [15:0] and_240__out;
  coreir_and #(.width(16)) and_240(
    .in0(and_240__in0),
    .in1(and_240__in1),
    .out(and_240__out)
  );

  //Wire declarations for instance 'and_242' (Module coreir_and)
  wire [15:0] and_242__in0;
  wire [15:0] and_242__in1;
  wire [15:0] and_242__out;
  coreir_and #(.width(16)) and_242(
    .in0(and_242__in0),
    .in1(and_242__in1),
    .out(and_242__out)
  );

  //Wire declarations for instance 'and_244' (Module coreir_and)
  wire [15:0] and_244__in0;
  wire [15:0] and_244__in1;
  wire [15:0] and_244__out;
  coreir_and #(.width(16)) and_244(
    .in0(and_244__in0),
    .in1(and_244__in1),
    .out(and_244__out)
  );

  //Wire declarations for instance 'and_246' (Module coreir_and)
  wire [15:0] and_246__in0;
  wire [15:0] and_246__in1;
  wire [15:0] and_246__out;
  coreir_and #(.width(16)) and_246(
    .in0(and_246__in0),
    .in1(and_246__in1),
    .out(and_246__out)
  );

  //Wire declarations for instance 'and_248' (Module coreir_and)
  wire [15:0] and_248__in0;
  wire [15:0] and_248__in1;
  wire [15:0] and_248__out;
  coreir_and #(.width(16)) and_248(
    .in0(and_248__in0),
    .in1(and_248__in1),
    .out(and_248__out)
  );

  //Wire declarations for instance 'and_250' (Module coreir_and)
  wire [15:0] and_250__in0;
  wire [15:0] and_250__in1;
  wire [15:0] and_250__out;
  coreir_and #(.width(16)) and_250(
    .in0(and_250__in0),
    .in1(and_250__in1),
    .out(and_250__out)
  );

  //Wire declarations for instance 'and_252' (Module coreir_and)
  wire [15:0] and_252__in0;
  wire [15:0] and_252__in1;
  wire [15:0] and_252__out;
  coreir_and #(.width(16)) and_252(
    .in0(and_252__in0),
    .in1(and_252__in1),
    .out(and_252__out)
  );

  //Wire declarations for instance 'and_254' (Module coreir_and)
  wire [15:0] and_254__in0;
  wire [15:0] and_254__in1;
  wire [15:0] and_254__out;
  coreir_and #(.width(16)) and_254(
    .in0(and_254__in0),
    .in1(and_254__in1),
    .out(and_254__out)
  );

  //Wire declarations for instance 'and_256' (Module coreir_and)
  wire [15:0] and_256__in0;
  wire [15:0] and_256__in1;
  wire [15:0] and_256__out;
  coreir_and #(.width(16)) and_256(
    .in0(and_256__in0),
    .in1(and_256__in1),
    .out(and_256__out)
  );

  //Wire declarations for instance 'and_258' (Module coreir_and)
  wire [15:0] and_258__in0;
  wire [15:0] and_258__in1;
  wire [15:0] and_258__out;
  coreir_and #(.width(16)) and_258(
    .in0(and_258__in0),
    .in1(and_258__in1),
    .out(and_258__out)
  );

  //Wire declarations for instance 'and_26' (Module coreir_and)
  wire [15:0] and_26__in0;
  wire [15:0] and_26__in1;
  wire [15:0] and_26__out;
  coreir_and #(.width(16)) and_26(
    .in0(and_26__in0),
    .in1(and_26__in1),
    .out(and_26__out)
  );

  //Wire declarations for instance 'and_260' (Module coreir_and)
  wire [15:0] and_260__in0;
  wire [15:0] and_260__in1;
  wire [15:0] and_260__out;
  coreir_and #(.width(16)) and_260(
    .in0(and_260__in0),
    .in1(and_260__in1),
    .out(and_260__out)
  );

  //Wire declarations for instance 'and_262' (Module coreir_and)
  wire [15:0] and_262__in0;
  wire [15:0] and_262__in1;
  wire [15:0] and_262__out;
  coreir_and #(.width(16)) and_262(
    .in0(and_262__in0),
    .in1(and_262__in1),
    .out(and_262__out)
  );

  //Wire declarations for instance 'and_264' (Module coreir_and)
  wire [15:0] and_264__in0;
  wire [15:0] and_264__in1;
  wire [15:0] and_264__out;
  coreir_and #(.width(16)) and_264(
    .in0(and_264__in0),
    .in1(and_264__in1),
    .out(and_264__out)
  );

  //Wire declarations for instance 'and_266' (Module coreir_and)
  wire [15:0] and_266__in0;
  wire [15:0] and_266__in1;
  wire [15:0] and_266__out;
  coreir_and #(.width(16)) and_266(
    .in0(and_266__in0),
    .in1(and_266__in1),
    .out(and_266__out)
  );

  //Wire declarations for instance 'and_268' (Module coreir_and)
  wire [15:0] and_268__in0;
  wire [15:0] and_268__in1;
  wire [15:0] and_268__out;
  coreir_and #(.width(16)) and_268(
    .in0(and_268__in0),
    .in1(and_268__in1),
    .out(and_268__out)
  );

  //Wire declarations for instance 'and_270' (Module coreir_and)
  wire [15:0] and_270__in0;
  wire [15:0] and_270__in1;
  wire [15:0] and_270__out;
  coreir_and #(.width(16)) and_270(
    .in0(and_270__in0),
    .in1(and_270__in1),
    .out(and_270__out)
  );

  //Wire declarations for instance 'and_272' (Module coreir_and)
  wire [15:0] and_272__in0;
  wire [15:0] and_272__in1;
  wire [15:0] and_272__out;
  coreir_and #(.width(16)) and_272(
    .in0(and_272__in0),
    .in1(and_272__in1),
    .out(and_272__out)
  );

  //Wire declarations for instance 'and_274' (Module coreir_and)
  wire [15:0] and_274__in0;
  wire [15:0] and_274__in1;
  wire [15:0] and_274__out;
  coreir_and #(.width(16)) and_274(
    .in0(and_274__in0),
    .in1(and_274__in1),
    .out(and_274__out)
  );

  //Wire declarations for instance 'and_276' (Module coreir_and)
  wire [15:0] and_276__in0;
  wire [15:0] and_276__in1;
  wire [15:0] and_276__out;
  coreir_and #(.width(16)) and_276(
    .in0(and_276__in0),
    .in1(and_276__in1),
    .out(and_276__out)
  );

  //Wire declarations for instance 'and_278' (Module coreir_and)
  wire [15:0] and_278__in0;
  wire [15:0] and_278__in1;
  wire [15:0] and_278__out;
  coreir_and #(.width(16)) and_278(
    .in0(and_278__in0),
    .in1(and_278__in1),
    .out(and_278__out)
  );

  //Wire declarations for instance 'and_28' (Module coreir_and)
  wire [15:0] and_28__in0;
  wire [15:0] and_28__in1;
  wire [15:0] and_28__out;
  coreir_and #(.width(16)) and_28(
    .in0(and_28__in0),
    .in1(and_28__in1),
    .out(and_28__out)
  );

  //Wire declarations for instance 'and_280' (Module coreir_and)
  wire [15:0] and_280__in0;
  wire [15:0] and_280__in1;
  wire [15:0] and_280__out;
  coreir_and #(.width(16)) and_280(
    .in0(and_280__in0),
    .in1(and_280__in1),
    .out(and_280__out)
  );

  //Wire declarations for instance 'and_282' (Module coreir_and)
  wire [15:0] and_282__in0;
  wire [15:0] and_282__in1;
  wire [15:0] and_282__out;
  coreir_and #(.width(16)) and_282(
    .in0(and_282__in0),
    .in1(and_282__in1),
    .out(and_282__out)
  );

  //Wire declarations for instance 'and_284' (Module coreir_and)
  wire [15:0] and_284__in0;
  wire [15:0] and_284__in1;
  wire [15:0] and_284__out;
  coreir_and #(.width(16)) and_284(
    .in0(and_284__in0),
    .in1(and_284__in1),
    .out(and_284__out)
  );

  //Wire declarations for instance 'and_286' (Module coreir_and)
  wire [15:0] and_286__in0;
  wire [15:0] and_286__in1;
  wire [15:0] and_286__out;
  coreir_and #(.width(16)) and_286(
    .in0(and_286__in0),
    .in1(and_286__in1),
    .out(and_286__out)
  );

  //Wire declarations for instance 'and_288' (Module coreir_and)
  wire [15:0] and_288__in0;
  wire [15:0] and_288__in1;
  wire [15:0] and_288__out;
  coreir_and #(.width(16)) and_288(
    .in0(and_288__in0),
    .in1(and_288__in1),
    .out(and_288__out)
  );

  //Wire declarations for instance 'and_290' (Module coreir_and)
  wire [15:0] and_290__in0;
  wire [15:0] and_290__in1;
  wire [15:0] and_290__out;
  coreir_and #(.width(16)) and_290(
    .in0(and_290__in0),
    .in1(and_290__in1),
    .out(and_290__out)
  );

  //Wire declarations for instance 'and_292' (Module coreir_and)
  wire [15:0] and_292__in0;
  wire [15:0] and_292__in1;
  wire [15:0] and_292__out;
  coreir_and #(.width(16)) and_292(
    .in0(and_292__in0),
    .in1(and_292__in1),
    .out(and_292__out)
  );

  //Wire declarations for instance 'and_294' (Module coreir_and)
  wire [15:0] and_294__in0;
  wire [15:0] and_294__in1;
  wire [15:0] and_294__out;
  coreir_and #(.width(16)) and_294(
    .in0(and_294__in0),
    .in1(and_294__in1),
    .out(and_294__out)
  );

  //Wire declarations for instance 'and_296' (Module coreir_and)
  wire [15:0] and_296__in0;
  wire [15:0] and_296__in1;
  wire [15:0] and_296__out;
  coreir_and #(.width(16)) and_296(
    .in0(and_296__in0),
    .in1(and_296__in1),
    .out(and_296__out)
  );

  //Wire declarations for instance 'and_298' (Module coreir_and)
  wire [15:0] and_298__in0;
  wire [15:0] and_298__in1;
  wire [15:0] and_298__out;
  coreir_and #(.width(16)) and_298(
    .in0(and_298__in0),
    .in1(and_298__in1),
    .out(and_298__out)
  );

  //Wire declarations for instance 'and_30' (Module coreir_and)
  wire [15:0] and_30__in0;
  wire [15:0] and_30__in1;
  wire [15:0] and_30__out;
  coreir_and #(.width(16)) and_30(
    .in0(and_30__in0),
    .in1(and_30__in1),
    .out(and_30__out)
  );

  //Wire declarations for instance 'and_300' (Module coreir_and)
  wire [15:0] and_300__in0;
  wire [15:0] and_300__in1;
  wire [15:0] and_300__out;
  coreir_and #(.width(16)) and_300(
    .in0(and_300__in0),
    .in1(and_300__in1),
    .out(and_300__out)
  );

  //Wire declarations for instance 'and_302' (Module coreir_and)
  wire [15:0] and_302__in0;
  wire [15:0] and_302__in1;
  wire [15:0] and_302__out;
  coreir_and #(.width(16)) and_302(
    .in0(and_302__in0),
    .in1(and_302__in1),
    .out(and_302__out)
  );

  //Wire declarations for instance 'and_304' (Module coreir_and)
  wire [15:0] and_304__in0;
  wire [15:0] and_304__in1;
  wire [15:0] and_304__out;
  coreir_and #(.width(16)) and_304(
    .in0(and_304__in0),
    .in1(and_304__in1),
    .out(and_304__out)
  );

  //Wire declarations for instance 'and_306' (Module coreir_and)
  wire [15:0] and_306__in0;
  wire [15:0] and_306__in1;
  wire [15:0] and_306__out;
  coreir_and #(.width(16)) and_306(
    .in0(and_306__in0),
    .in1(and_306__in1),
    .out(and_306__out)
  );

  //Wire declarations for instance 'and_308' (Module coreir_and)
  wire [15:0] and_308__in0;
  wire [15:0] and_308__in1;
  wire [15:0] and_308__out;
  coreir_and #(.width(16)) and_308(
    .in0(and_308__in0),
    .in1(and_308__in1),
    .out(and_308__out)
  );

  //Wire declarations for instance 'and_310' (Module coreir_and)
  wire [15:0] and_310__in0;
  wire [15:0] and_310__in1;
  wire [15:0] and_310__out;
  coreir_and #(.width(16)) and_310(
    .in0(and_310__in0),
    .in1(and_310__in1),
    .out(and_310__out)
  );

  //Wire declarations for instance 'and_312' (Module coreir_and)
  wire [15:0] and_312__in0;
  wire [15:0] and_312__in1;
  wire [15:0] and_312__out;
  coreir_and #(.width(16)) and_312(
    .in0(and_312__in0),
    .in1(and_312__in1),
    .out(and_312__out)
  );

  //Wire declarations for instance 'and_314' (Module coreir_and)
  wire [15:0] and_314__in0;
  wire [15:0] and_314__in1;
  wire [15:0] and_314__out;
  coreir_and #(.width(16)) and_314(
    .in0(and_314__in0),
    .in1(and_314__in1),
    .out(and_314__out)
  );

  //Wire declarations for instance 'and_316' (Module coreir_and)
  wire [15:0] and_316__in0;
  wire [15:0] and_316__in1;
  wire [15:0] and_316__out;
  coreir_and #(.width(16)) and_316(
    .in0(and_316__in0),
    .in1(and_316__in1),
    .out(and_316__out)
  );

  //Wire declarations for instance 'and_318' (Module coreir_and)
  wire [15:0] and_318__in0;
  wire [15:0] and_318__in1;
  wire [15:0] and_318__out;
  coreir_and #(.width(16)) and_318(
    .in0(and_318__in0),
    .in1(and_318__in1),
    .out(and_318__out)
  );

  //Wire declarations for instance 'and_32' (Module coreir_and)
  wire [15:0] and_32__in0;
  wire [15:0] and_32__in1;
  wire [15:0] and_32__out;
  coreir_and #(.width(16)) and_32(
    .in0(and_32__in0),
    .in1(and_32__in1),
    .out(and_32__out)
  );

  //Wire declarations for instance 'and_320' (Module coreir_and)
  wire [15:0] and_320__in0;
  wire [15:0] and_320__in1;
  wire [15:0] and_320__out;
  coreir_and #(.width(16)) and_320(
    .in0(and_320__in0),
    .in1(and_320__in1),
    .out(and_320__out)
  );

  //Wire declarations for instance 'and_322' (Module coreir_and)
  wire [15:0] and_322__in0;
  wire [15:0] and_322__in1;
  wire [15:0] and_322__out;
  coreir_and #(.width(16)) and_322(
    .in0(and_322__in0),
    .in1(and_322__in1),
    .out(and_322__out)
  );

  //Wire declarations for instance 'and_324' (Module coreir_and)
  wire [15:0] and_324__in0;
  wire [15:0] and_324__in1;
  wire [15:0] and_324__out;
  coreir_and #(.width(16)) and_324(
    .in0(and_324__in0),
    .in1(and_324__in1),
    .out(and_324__out)
  );

  //Wire declarations for instance 'and_326' (Module coreir_and)
  wire [15:0] and_326__in0;
  wire [15:0] and_326__in1;
  wire [15:0] and_326__out;
  coreir_and #(.width(16)) and_326(
    .in0(and_326__in0),
    .in1(and_326__in1),
    .out(and_326__out)
  );

  //Wire declarations for instance 'and_328' (Module coreir_and)
  wire [15:0] and_328__in0;
  wire [15:0] and_328__in1;
  wire [15:0] and_328__out;
  coreir_and #(.width(16)) and_328(
    .in0(and_328__in0),
    .in1(and_328__in1),
    .out(and_328__out)
  );

  //Wire declarations for instance 'and_330' (Module coreir_and)
  wire [15:0] and_330__in0;
  wire [15:0] and_330__in1;
  wire [15:0] and_330__out;
  coreir_and #(.width(16)) and_330(
    .in0(and_330__in0),
    .in1(and_330__in1),
    .out(and_330__out)
  );

  //Wire declarations for instance 'and_332' (Module coreir_and)
  wire [15:0] and_332__in0;
  wire [15:0] and_332__in1;
  wire [15:0] and_332__out;
  coreir_and #(.width(16)) and_332(
    .in0(and_332__in0),
    .in1(and_332__in1),
    .out(and_332__out)
  );

  //Wire declarations for instance 'and_334' (Module coreir_and)
  wire [15:0] and_334__in0;
  wire [15:0] and_334__in1;
  wire [15:0] and_334__out;
  coreir_and #(.width(16)) and_334(
    .in0(and_334__in0),
    .in1(and_334__in1),
    .out(and_334__out)
  );

  //Wire declarations for instance 'and_336' (Module coreir_and)
  wire [15:0] and_336__in0;
  wire [15:0] and_336__in1;
  wire [15:0] and_336__out;
  coreir_and #(.width(16)) and_336(
    .in0(and_336__in0),
    .in1(and_336__in1),
    .out(and_336__out)
  );

  //Wire declarations for instance 'and_338' (Module coreir_and)
  wire [15:0] and_338__in0;
  wire [15:0] and_338__in1;
  wire [15:0] and_338__out;
  coreir_and #(.width(16)) and_338(
    .in0(and_338__in0),
    .in1(and_338__in1),
    .out(and_338__out)
  );

  //Wire declarations for instance 'and_34' (Module coreir_and)
  wire [15:0] and_34__in0;
  wire [15:0] and_34__in1;
  wire [15:0] and_34__out;
  coreir_and #(.width(16)) and_34(
    .in0(and_34__in0),
    .in1(and_34__in1),
    .out(and_34__out)
  );

  //Wire declarations for instance 'and_340' (Module coreir_and)
  wire [15:0] and_340__in0;
  wire [15:0] and_340__in1;
  wire [15:0] and_340__out;
  coreir_and #(.width(16)) and_340(
    .in0(and_340__in0),
    .in1(and_340__in1),
    .out(and_340__out)
  );

  //Wire declarations for instance 'and_342' (Module coreir_and)
  wire [15:0] and_342__in0;
  wire [15:0] and_342__in1;
  wire [15:0] and_342__out;
  coreir_and #(.width(16)) and_342(
    .in0(and_342__in0),
    .in1(and_342__in1),
    .out(and_342__out)
  );

  //Wire declarations for instance 'and_344' (Module coreir_and)
  wire [15:0] and_344__in0;
  wire [15:0] and_344__in1;
  wire [15:0] and_344__out;
  coreir_and #(.width(16)) and_344(
    .in0(and_344__in0),
    .in1(and_344__in1),
    .out(and_344__out)
  );

  //Wire declarations for instance 'and_346' (Module coreir_and)
  wire [15:0] and_346__in0;
  wire [15:0] and_346__in1;
  wire [15:0] and_346__out;
  coreir_and #(.width(16)) and_346(
    .in0(and_346__in0),
    .in1(and_346__in1),
    .out(and_346__out)
  );

  //Wire declarations for instance 'and_348' (Module coreir_and)
  wire [15:0] and_348__in0;
  wire [15:0] and_348__in1;
  wire [15:0] and_348__out;
  coreir_and #(.width(16)) and_348(
    .in0(and_348__in0),
    .in1(and_348__in1),
    .out(and_348__out)
  );

  //Wire declarations for instance 'and_350' (Module coreir_and)
  wire [15:0] and_350__in0;
  wire [15:0] and_350__in1;
  wire [15:0] and_350__out;
  coreir_and #(.width(16)) and_350(
    .in0(and_350__in0),
    .in1(and_350__in1),
    .out(and_350__out)
  );

  //Wire declarations for instance 'and_352' (Module coreir_and)
  wire [15:0] and_352__in0;
  wire [15:0] and_352__in1;
  wire [15:0] and_352__out;
  coreir_and #(.width(16)) and_352(
    .in0(and_352__in0),
    .in1(and_352__in1),
    .out(and_352__out)
  );

  //Wire declarations for instance 'and_354' (Module coreir_and)
  wire [15:0] and_354__in0;
  wire [15:0] and_354__in1;
  wire [15:0] and_354__out;
  coreir_and #(.width(16)) and_354(
    .in0(and_354__in0),
    .in1(and_354__in1),
    .out(and_354__out)
  );

  //Wire declarations for instance 'and_356' (Module coreir_and)
  wire [15:0] and_356__in0;
  wire [15:0] and_356__in1;
  wire [15:0] and_356__out;
  coreir_and #(.width(16)) and_356(
    .in0(and_356__in0),
    .in1(and_356__in1),
    .out(and_356__out)
  );

  //Wire declarations for instance 'and_358' (Module coreir_and)
  wire [15:0] and_358__in0;
  wire [15:0] and_358__in1;
  wire [15:0] and_358__out;
  coreir_and #(.width(16)) and_358(
    .in0(and_358__in0),
    .in1(and_358__in1),
    .out(and_358__out)
  );

  //Wire declarations for instance 'and_36' (Module coreir_and)
  wire [15:0] and_36__in0;
  wire [15:0] and_36__in1;
  wire [15:0] and_36__out;
  coreir_and #(.width(16)) and_36(
    .in0(and_36__in0),
    .in1(and_36__in1),
    .out(and_36__out)
  );

  //Wire declarations for instance 'and_360' (Module coreir_and)
  wire [15:0] and_360__in0;
  wire [15:0] and_360__in1;
  wire [15:0] and_360__out;
  coreir_and #(.width(16)) and_360(
    .in0(and_360__in0),
    .in1(and_360__in1),
    .out(and_360__out)
  );

  //Wire declarations for instance 'and_362' (Module coreir_and)
  wire [15:0] and_362__in0;
  wire [15:0] and_362__in1;
  wire [15:0] and_362__out;
  coreir_and #(.width(16)) and_362(
    .in0(and_362__in0),
    .in1(and_362__in1),
    .out(and_362__out)
  );

  //Wire declarations for instance 'and_364' (Module coreir_and)
  wire [15:0] and_364__in0;
  wire [15:0] and_364__in1;
  wire [15:0] and_364__out;
  coreir_and #(.width(16)) and_364(
    .in0(and_364__in0),
    .in1(and_364__in1),
    .out(and_364__out)
  );

  //Wire declarations for instance 'and_366' (Module coreir_and)
  wire [15:0] and_366__in0;
  wire [15:0] and_366__in1;
  wire [15:0] and_366__out;
  coreir_and #(.width(16)) and_366(
    .in0(and_366__in0),
    .in1(and_366__in1),
    .out(and_366__out)
  );

  //Wire declarations for instance 'and_368' (Module coreir_and)
  wire [15:0] and_368__in0;
  wire [15:0] and_368__in1;
  wire [15:0] and_368__out;
  coreir_and #(.width(16)) and_368(
    .in0(and_368__in0),
    .in1(and_368__in1),
    .out(and_368__out)
  );

  //Wire declarations for instance 'and_370' (Module coreir_and)
  wire [15:0] and_370__in0;
  wire [15:0] and_370__in1;
  wire [15:0] and_370__out;
  coreir_and #(.width(16)) and_370(
    .in0(and_370__in0),
    .in1(and_370__in1),
    .out(and_370__out)
  );

  //Wire declarations for instance 'and_372' (Module coreir_and)
  wire [15:0] and_372__in0;
  wire [15:0] and_372__in1;
  wire [15:0] and_372__out;
  coreir_and #(.width(16)) and_372(
    .in0(and_372__in0),
    .in1(and_372__in1),
    .out(and_372__out)
  );

  //Wire declarations for instance 'and_374' (Module coreir_and)
  wire [15:0] and_374__in0;
  wire [15:0] and_374__in1;
  wire [15:0] and_374__out;
  coreir_and #(.width(16)) and_374(
    .in0(and_374__in0),
    .in1(and_374__in1),
    .out(and_374__out)
  );

  //Wire declarations for instance 'and_376' (Module coreir_and)
  wire [15:0] and_376__in0;
  wire [15:0] and_376__in1;
  wire [15:0] and_376__out;
  coreir_and #(.width(16)) and_376(
    .in0(and_376__in0),
    .in1(and_376__in1),
    .out(and_376__out)
  );

  //Wire declarations for instance 'and_378' (Module coreir_and)
  wire [15:0] and_378__in0;
  wire [15:0] and_378__in1;
  wire [15:0] and_378__out;
  coreir_and #(.width(16)) and_378(
    .in0(and_378__in0),
    .in1(and_378__in1),
    .out(and_378__out)
  );

  //Wire declarations for instance 'and_38' (Module coreir_and)
  wire [15:0] and_38__in0;
  wire [15:0] and_38__in1;
  wire [15:0] and_38__out;
  coreir_and #(.width(16)) and_38(
    .in0(and_38__in0),
    .in1(and_38__in1),
    .out(and_38__out)
  );

  //Wire declarations for instance 'and_380' (Module coreir_and)
  wire [15:0] and_380__in0;
  wire [15:0] and_380__in1;
  wire [15:0] and_380__out;
  coreir_and #(.width(16)) and_380(
    .in0(and_380__in0),
    .in1(and_380__in1),
    .out(and_380__out)
  );

  //Wire declarations for instance 'and_382' (Module coreir_and)
  wire [15:0] and_382__in0;
  wire [15:0] and_382__in1;
  wire [15:0] and_382__out;
  coreir_and #(.width(16)) and_382(
    .in0(and_382__in0),
    .in1(and_382__in1),
    .out(and_382__out)
  );

  //Wire declarations for instance 'and_384' (Module coreir_and)
  wire [15:0] and_384__in0;
  wire [15:0] and_384__in1;
  wire [15:0] and_384__out;
  coreir_and #(.width(16)) and_384(
    .in0(and_384__in0),
    .in1(and_384__in1),
    .out(and_384__out)
  );

  //Wire declarations for instance 'and_386' (Module coreir_and)
  wire [15:0] and_386__in0;
  wire [15:0] and_386__in1;
  wire [15:0] and_386__out;
  coreir_and #(.width(16)) and_386(
    .in0(and_386__in0),
    .in1(and_386__in1),
    .out(and_386__out)
  );

  //Wire declarations for instance 'and_388' (Module coreir_and)
  wire [15:0] and_388__in0;
  wire [15:0] and_388__in1;
  wire [15:0] and_388__out;
  coreir_and #(.width(16)) and_388(
    .in0(and_388__in0),
    .in1(and_388__in1),
    .out(and_388__out)
  );

  //Wire declarations for instance 'and_390' (Module coreir_and)
  wire [15:0] and_390__in0;
  wire [15:0] and_390__in1;
  wire [15:0] and_390__out;
  coreir_and #(.width(16)) and_390(
    .in0(and_390__in0),
    .in1(and_390__in1),
    .out(and_390__out)
  );

  //Wire declarations for instance 'and_392' (Module coreir_and)
  wire [15:0] and_392__in0;
  wire [15:0] and_392__in1;
  wire [15:0] and_392__out;
  coreir_and #(.width(16)) and_392(
    .in0(and_392__in0),
    .in1(and_392__in1),
    .out(and_392__out)
  );

  //Wire declarations for instance 'and_394' (Module coreir_and)
  wire [15:0] and_394__in0;
  wire [15:0] and_394__in1;
  wire [15:0] and_394__out;
  coreir_and #(.width(16)) and_394(
    .in0(and_394__in0),
    .in1(and_394__in1),
    .out(and_394__out)
  );

  //Wire declarations for instance 'and_396' (Module coreir_and)
  wire [15:0] and_396__in0;
  wire [15:0] and_396__in1;
  wire [15:0] and_396__out;
  coreir_and #(.width(16)) and_396(
    .in0(and_396__in0),
    .in1(and_396__in1),
    .out(and_396__out)
  );

  //Wire declarations for instance 'and_398' (Module coreir_and)
  wire [15:0] and_398__in0;
  wire [15:0] and_398__in1;
  wire [15:0] and_398__out;
  coreir_and #(.width(16)) and_398(
    .in0(and_398__in0),
    .in1(and_398__in1),
    .out(and_398__out)
  );

  //Wire declarations for instance 'and_4' (Module coreir_and)
  wire [15:0] and_4__in0;
  wire [15:0] and_4__in1;
  wire [15:0] and_4__out;
  coreir_and #(.width(16)) and_4(
    .in0(and_4__in0),
    .in1(and_4__in1),
    .out(and_4__out)
  );

  //Wire declarations for instance 'and_40' (Module coreir_and)
  wire [15:0] and_40__in0;
  wire [15:0] and_40__in1;
  wire [15:0] and_40__out;
  coreir_and #(.width(16)) and_40(
    .in0(and_40__in0),
    .in1(and_40__in1),
    .out(and_40__out)
  );

  //Wire declarations for instance 'and_400' (Module coreir_and)
  wire [15:0] and_400__in0;
  wire [15:0] and_400__in1;
  wire [15:0] and_400__out;
  coreir_and #(.width(16)) and_400(
    .in0(and_400__in0),
    .in1(and_400__in1),
    .out(and_400__out)
  );

  //Wire declarations for instance 'and_402' (Module coreir_and)
  wire [15:0] and_402__in0;
  wire [15:0] and_402__in1;
  wire [15:0] and_402__out;
  coreir_and #(.width(16)) and_402(
    .in0(and_402__in0),
    .in1(and_402__in1),
    .out(and_402__out)
  );

  //Wire declarations for instance 'and_404' (Module coreir_and)
  wire [15:0] and_404__in0;
  wire [15:0] and_404__in1;
  wire [15:0] and_404__out;
  coreir_and #(.width(16)) and_404(
    .in0(and_404__in0),
    .in1(and_404__in1),
    .out(and_404__out)
  );

  //Wire declarations for instance 'and_406' (Module coreir_and)
  wire [15:0] and_406__in0;
  wire [15:0] and_406__in1;
  wire [15:0] and_406__out;
  coreir_and #(.width(16)) and_406(
    .in0(and_406__in0),
    .in1(and_406__in1),
    .out(and_406__out)
  );

  //Wire declarations for instance 'and_408' (Module coreir_and)
  wire [15:0] and_408__in0;
  wire [15:0] and_408__in1;
  wire [15:0] and_408__out;
  coreir_and #(.width(16)) and_408(
    .in0(and_408__in0),
    .in1(and_408__in1),
    .out(and_408__out)
  );

  //Wire declarations for instance 'and_410' (Module coreir_and)
  wire [15:0] and_410__in0;
  wire [15:0] and_410__in1;
  wire [15:0] and_410__out;
  coreir_and #(.width(16)) and_410(
    .in0(and_410__in0),
    .in1(and_410__in1),
    .out(and_410__out)
  );

  //Wire declarations for instance 'and_412' (Module coreir_and)
  wire [15:0] and_412__in0;
  wire [15:0] and_412__in1;
  wire [15:0] and_412__out;
  coreir_and #(.width(16)) and_412(
    .in0(and_412__in0),
    .in1(and_412__in1),
    .out(and_412__out)
  );

  //Wire declarations for instance 'and_414' (Module coreir_and)
  wire [15:0] and_414__in0;
  wire [15:0] and_414__in1;
  wire [15:0] and_414__out;
  coreir_and #(.width(16)) and_414(
    .in0(and_414__in0),
    .in1(and_414__in1),
    .out(and_414__out)
  );

  //Wire declarations for instance 'and_416' (Module coreir_and)
  wire [15:0] and_416__in0;
  wire [15:0] and_416__in1;
  wire [15:0] and_416__out;
  coreir_and #(.width(16)) and_416(
    .in0(and_416__in0),
    .in1(and_416__in1),
    .out(and_416__out)
  );

  //Wire declarations for instance 'and_418' (Module coreir_and)
  wire [15:0] and_418__in0;
  wire [15:0] and_418__in1;
  wire [15:0] and_418__out;
  coreir_and #(.width(16)) and_418(
    .in0(and_418__in0),
    .in1(and_418__in1),
    .out(and_418__out)
  );

  //Wire declarations for instance 'and_42' (Module coreir_and)
  wire [15:0] and_42__in0;
  wire [15:0] and_42__in1;
  wire [15:0] and_42__out;
  coreir_and #(.width(16)) and_42(
    .in0(and_42__in0),
    .in1(and_42__in1),
    .out(and_42__out)
  );

  //Wire declarations for instance 'and_420' (Module coreir_and)
  wire [15:0] and_420__in0;
  wire [15:0] and_420__in1;
  wire [15:0] and_420__out;
  coreir_and #(.width(16)) and_420(
    .in0(and_420__in0),
    .in1(and_420__in1),
    .out(and_420__out)
  );

  //Wire declarations for instance 'and_422' (Module coreir_and)
  wire [15:0] and_422__in0;
  wire [15:0] and_422__in1;
  wire [15:0] and_422__out;
  coreir_and #(.width(16)) and_422(
    .in0(and_422__in0),
    .in1(and_422__in1),
    .out(and_422__out)
  );

  //Wire declarations for instance 'and_424' (Module coreir_and)
  wire [15:0] and_424__in0;
  wire [15:0] and_424__in1;
  wire [15:0] and_424__out;
  coreir_and #(.width(16)) and_424(
    .in0(and_424__in0),
    .in1(and_424__in1),
    .out(and_424__out)
  );

  //Wire declarations for instance 'and_426' (Module coreir_and)
  wire [15:0] and_426__in0;
  wire [15:0] and_426__in1;
  wire [15:0] and_426__out;
  coreir_and #(.width(16)) and_426(
    .in0(and_426__in0),
    .in1(and_426__in1),
    .out(and_426__out)
  );

  //Wire declarations for instance 'and_428' (Module coreir_and)
  wire [15:0] and_428__in0;
  wire [15:0] and_428__in1;
  wire [15:0] and_428__out;
  coreir_and #(.width(16)) and_428(
    .in0(and_428__in0),
    .in1(and_428__in1),
    .out(and_428__out)
  );

  //Wire declarations for instance 'and_430' (Module coreir_and)
  wire [15:0] and_430__in0;
  wire [15:0] and_430__in1;
  wire [15:0] and_430__out;
  coreir_and #(.width(16)) and_430(
    .in0(and_430__in0),
    .in1(and_430__in1),
    .out(and_430__out)
  );

  //Wire declarations for instance 'and_432' (Module coreir_and)
  wire [15:0] and_432__in0;
  wire [15:0] and_432__in1;
  wire [15:0] and_432__out;
  coreir_and #(.width(16)) and_432(
    .in0(and_432__in0),
    .in1(and_432__in1),
    .out(and_432__out)
  );

  //Wire declarations for instance 'and_434' (Module coreir_and)
  wire [15:0] and_434__in0;
  wire [15:0] and_434__in1;
  wire [15:0] and_434__out;
  coreir_and #(.width(16)) and_434(
    .in0(and_434__in0),
    .in1(and_434__in1),
    .out(and_434__out)
  );

  //Wire declarations for instance 'and_436' (Module coreir_and)
  wire [15:0] and_436__in0;
  wire [15:0] and_436__in1;
  wire [15:0] and_436__out;
  coreir_and #(.width(16)) and_436(
    .in0(and_436__in0),
    .in1(and_436__in1),
    .out(and_436__out)
  );

  //Wire declarations for instance 'and_438' (Module coreir_and)
  wire [15:0] and_438__in0;
  wire [15:0] and_438__in1;
  wire [15:0] and_438__out;
  coreir_and #(.width(16)) and_438(
    .in0(and_438__in0),
    .in1(and_438__in1),
    .out(and_438__out)
  );

  //Wire declarations for instance 'and_44' (Module coreir_and)
  wire [15:0] and_44__in0;
  wire [15:0] and_44__in1;
  wire [15:0] and_44__out;
  coreir_and #(.width(16)) and_44(
    .in0(and_44__in0),
    .in1(and_44__in1),
    .out(and_44__out)
  );

  //Wire declarations for instance 'and_440' (Module coreir_and)
  wire [15:0] and_440__in0;
  wire [15:0] and_440__in1;
  wire [15:0] and_440__out;
  coreir_and #(.width(16)) and_440(
    .in0(and_440__in0),
    .in1(and_440__in1),
    .out(and_440__out)
  );

  //Wire declarations for instance 'and_442' (Module coreir_and)
  wire [15:0] and_442__in0;
  wire [15:0] and_442__in1;
  wire [15:0] and_442__out;
  coreir_and #(.width(16)) and_442(
    .in0(and_442__in0),
    .in1(and_442__in1),
    .out(and_442__out)
  );

  //Wire declarations for instance 'and_444' (Module coreir_and)
  wire [15:0] and_444__in0;
  wire [15:0] and_444__in1;
  wire [15:0] and_444__out;
  coreir_and #(.width(16)) and_444(
    .in0(and_444__in0),
    .in1(and_444__in1),
    .out(and_444__out)
  );

  //Wire declarations for instance 'and_446' (Module coreir_and)
  wire [15:0] and_446__in0;
  wire [15:0] and_446__in1;
  wire [15:0] and_446__out;
  coreir_and #(.width(16)) and_446(
    .in0(and_446__in0),
    .in1(and_446__in1),
    .out(and_446__out)
  );

  //Wire declarations for instance 'and_448' (Module coreir_and)
  wire [15:0] and_448__in0;
  wire [15:0] and_448__in1;
  wire [15:0] and_448__out;
  coreir_and #(.width(16)) and_448(
    .in0(and_448__in0),
    .in1(and_448__in1),
    .out(and_448__out)
  );

  //Wire declarations for instance 'and_450' (Module coreir_and)
  wire [15:0] and_450__in0;
  wire [15:0] and_450__in1;
  wire [15:0] and_450__out;
  coreir_and #(.width(16)) and_450(
    .in0(and_450__in0),
    .in1(and_450__in1),
    .out(and_450__out)
  );

  //Wire declarations for instance 'and_452' (Module coreir_and)
  wire [15:0] and_452__in0;
  wire [15:0] and_452__in1;
  wire [15:0] and_452__out;
  coreir_and #(.width(16)) and_452(
    .in0(and_452__in0),
    .in1(and_452__in1),
    .out(and_452__out)
  );

  //Wire declarations for instance 'and_454' (Module coreir_and)
  wire [15:0] and_454__in0;
  wire [15:0] and_454__in1;
  wire [15:0] and_454__out;
  coreir_and #(.width(16)) and_454(
    .in0(and_454__in0),
    .in1(and_454__in1),
    .out(and_454__out)
  );

  //Wire declarations for instance 'and_456' (Module coreir_and)
  wire [15:0] and_456__in0;
  wire [15:0] and_456__in1;
  wire [15:0] and_456__out;
  coreir_and #(.width(16)) and_456(
    .in0(and_456__in0),
    .in1(and_456__in1),
    .out(and_456__out)
  );

  //Wire declarations for instance 'and_458' (Module coreir_and)
  wire [15:0] and_458__in0;
  wire [15:0] and_458__in1;
  wire [15:0] and_458__out;
  coreir_and #(.width(16)) and_458(
    .in0(and_458__in0),
    .in1(and_458__in1),
    .out(and_458__out)
  );

  //Wire declarations for instance 'and_46' (Module coreir_and)
  wire [15:0] and_46__in0;
  wire [15:0] and_46__in1;
  wire [15:0] and_46__out;
  coreir_and #(.width(16)) and_46(
    .in0(and_46__in0),
    .in1(and_46__in1),
    .out(and_46__out)
  );

  //Wire declarations for instance 'and_460' (Module coreir_and)
  wire [15:0] and_460__in0;
  wire [15:0] and_460__in1;
  wire [15:0] and_460__out;
  coreir_and #(.width(16)) and_460(
    .in0(and_460__in0),
    .in1(and_460__in1),
    .out(and_460__out)
  );

  //Wire declarations for instance 'and_462' (Module coreir_and)
  wire [15:0] and_462__in0;
  wire [15:0] and_462__in1;
  wire [15:0] and_462__out;
  coreir_and #(.width(16)) and_462(
    .in0(and_462__in0),
    .in1(and_462__in1),
    .out(and_462__out)
  );

  //Wire declarations for instance 'and_464' (Module coreir_and)
  wire [15:0] and_464__in0;
  wire [15:0] and_464__in1;
  wire [15:0] and_464__out;
  coreir_and #(.width(16)) and_464(
    .in0(and_464__in0),
    .in1(and_464__in1),
    .out(and_464__out)
  );

  //Wire declarations for instance 'and_466' (Module coreir_and)
  wire [15:0] and_466__in0;
  wire [15:0] and_466__in1;
  wire [15:0] and_466__out;
  coreir_and #(.width(16)) and_466(
    .in0(and_466__in0),
    .in1(and_466__in1),
    .out(and_466__out)
  );

  //Wire declarations for instance 'and_468' (Module coreir_and)
  wire [15:0] and_468__in0;
  wire [15:0] and_468__in1;
  wire [15:0] and_468__out;
  coreir_and #(.width(16)) and_468(
    .in0(and_468__in0),
    .in1(and_468__in1),
    .out(and_468__out)
  );

  //Wire declarations for instance 'and_470' (Module coreir_and)
  wire [15:0] and_470__in0;
  wire [15:0] and_470__in1;
  wire [15:0] and_470__out;
  coreir_and #(.width(16)) and_470(
    .in0(and_470__in0),
    .in1(and_470__in1),
    .out(and_470__out)
  );

  //Wire declarations for instance 'and_472' (Module coreir_and)
  wire [15:0] and_472__in0;
  wire [15:0] and_472__in1;
  wire [15:0] and_472__out;
  coreir_and #(.width(16)) and_472(
    .in0(and_472__in0),
    .in1(and_472__in1),
    .out(and_472__out)
  );

  //Wire declarations for instance 'and_474' (Module coreir_and)
  wire [15:0] and_474__in0;
  wire [15:0] and_474__in1;
  wire [15:0] and_474__out;
  coreir_and #(.width(16)) and_474(
    .in0(and_474__in0),
    .in1(and_474__in1),
    .out(and_474__out)
  );

  //Wire declarations for instance 'and_476' (Module coreir_and)
  wire [15:0] and_476__in0;
  wire [15:0] and_476__in1;
  wire [15:0] and_476__out;
  coreir_and #(.width(16)) and_476(
    .in0(and_476__in0),
    .in1(and_476__in1),
    .out(and_476__out)
  );

  //Wire declarations for instance 'and_478' (Module coreir_and)
  wire [15:0] and_478__in0;
  wire [15:0] and_478__in1;
  wire [15:0] and_478__out;
  coreir_and #(.width(16)) and_478(
    .in0(and_478__in0),
    .in1(and_478__in1),
    .out(and_478__out)
  );

  //Wire declarations for instance 'and_48' (Module coreir_and)
  wire [15:0] and_48__in0;
  wire [15:0] and_48__in1;
  wire [15:0] and_48__out;
  coreir_and #(.width(16)) and_48(
    .in0(and_48__in0),
    .in1(and_48__in1),
    .out(and_48__out)
  );

  //Wire declarations for instance 'and_480' (Module coreir_and)
  wire [15:0] and_480__in0;
  wire [15:0] and_480__in1;
  wire [15:0] and_480__out;
  coreir_and #(.width(16)) and_480(
    .in0(and_480__in0),
    .in1(and_480__in1),
    .out(and_480__out)
  );

  //Wire declarations for instance 'and_482' (Module coreir_and)
  wire [15:0] and_482__in0;
  wire [15:0] and_482__in1;
  wire [15:0] and_482__out;
  coreir_and #(.width(16)) and_482(
    .in0(and_482__in0),
    .in1(and_482__in1),
    .out(and_482__out)
  );

  //Wire declarations for instance 'and_484' (Module coreir_and)
  wire [15:0] and_484__in0;
  wire [15:0] and_484__in1;
  wire [15:0] and_484__out;
  coreir_and #(.width(16)) and_484(
    .in0(and_484__in0),
    .in1(and_484__in1),
    .out(and_484__out)
  );

  //Wire declarations for instance 'and_486' (Module coreir_and)
  wire [15:0] and_486__in0;
  wire [15:0] and_486__in1;
  wire [15:0] and_486__out;
  coreir_and #(.width(16)) and_486(
    .in0(and_486__in0),
    .in1(and_486__in1),
    .out(and_486__out)
  );

  //Wire declarations for instance 'and_488' (Module coreir_and)
  wire [15:0] and_488__in0;
  wire [15:0] and_488__in1;
  wire [15:0] and_488__out;
  coreir_and #(.width(16)) and_488(
    .in0(and_488__in0),
    .in1(and_488__in1),
    .out(and_488__out)
  );

  //Wire declarations for instance 'and_490' (Module coreir_and)
  wire [15:0] and_490__in0;
  wire [15:0] and_490__in1;
  wire [15:0] and_490__out;
  coreir_and #(.width(16)) and_490(
    .in0(and_490__in0),
    .in1(and_490__in1),
    .out(and_490__out)
  );

  //Wire declarations for instance 'and_492' (Module coreir_and)
  wire [15:0] and_492__in0;
  wire [15:0] and_492__in1;
  wire [15:0] and_492__out;
  coreir_and #(.width(16)) and_492(
    .in0(and_492__in0),
    .in1(and_492__in1),
    .out(and_492__out)
  );

  //Wire declarations for instance 'and_494' (Module coreir_and)
  wire [15:0] and_494__in0;
  wire [15:0] and_494__in1;
  wire [15:0] and_494__out;
  coreir_and #(.width(16)) and_494(
    .in0(and_494__in0),
    .in1(and_494__in1),
    .out(and_494__out)
  );

  //Wire declarations for instance 'and_496' (Module coreir_and)
  wire [15:0] and_496__in0;
  wire [15:0] and_496__in1;
  wire [15:0] and_496__out;
  coreir_and #(.width(16)) and_496(
    .in0(and_496__in0),
    .in1(and_496__in1),
    .out(and_496__out)
  );

  //Wire declarations for instance 'and_498' (Module coreir_and)
  wire [15:0] and_498__in0;
  wire [15:0] and_498__in1;
  wire [15:0] and_498__out;
  coreir_and #(.width(16)) and_498(
    .in0(and_498__in0),
    .in1(and_498__in1),
    .out(and_498__out)
  );

  //Wire declarations for instance 'and_50' (Module coreir_and)
  wire [15:0] and_50__in0;
  wire [15:0] and_50__in1;
  wire [15:0] and_50__out;
  coreir_and #(.width(16)) and_50(
    .in0(and_50__in0),
    .in1(and_50__in1),
    .out(and_50__out)
  );

  //Wire declarations for instance 'and_500' (Module coreir_and)
  wire [15:0] and_500__in0;
  wire [15:0] and_500__in1;
  wire [15:0] and_500__out;
  coreir_and #(.width(16)) and_500(
    .in0(and_500__in0),
    .in1(and_500__in1),
    .out(and_500__out)
  );

  //Wire declarations for instance 'and_502' (Module coreir_and)
  wire [15:0] and_502__in0;
  wire [15:0] and_502__in1;
  wire [15:0] and_502__out;
  coreir_and #(.width(16)) and_502(
    .in0(and_502__in0),
    .in1(and_502__in1),
    .out(and_502__out)
  );

  //Wire declarations for instance 'and_504' (Module coreir_and)
  wire [15:0] and_504__in0;
  wire [15:0] and_504__in1;
  wire [15:0] and_504__out;
  coreir_and #(.width(16)) and_504(
    .in0(and_504__in0),
    .in1(and_504__in1),
    .out(and_504__out)
  );

  //Wire declarations for instance 'and_506' (Module coreir_and)
  wire [15:0] and_506__in0;
  wire [15:0] and_506__in1;
  wire [15:0] and_506__out;
  coreir_and #(.width(16)) and_506(
    .in0(and_506__in0),
    .in1(and_506__in1),
    .out(and_506__out)
  );

  //Wire declarations for instance 'and_508' (Module coreir_and)
  wire [15:0] and_508__in0;
  wire [15:0] and_508__in1;
  wire [15:0] and_508__out;
  coreir_and #(.width(16)) and_508(
    .in0(and_508__in0),
    .in1(and_508__in1),
    .out(and_508__out)
  );

  //Wire declarations for instance 'and_510' (Module coreir_and)
  wire [15:0] and_510__in0;
  wire [15:0] and_510__in1;
  wire [15:0] and_510__out;
  coreir_and #(.width(16)) and_510(
    .in0(and_510__in0),
    .in1(and_510__in1),
    .out(and_510__out)
  );

  //Wire declarations for instance 'and_512' (Module coreir_and)
  wire [15:0] and_512__in0;
  wire [15:0] and_512__in1;
  wire [15:0] and_512__out;
  coreir_and #(.width(16)) and_512(
    .in0(and_512__in0),
    .in1(and_512__in1),
    .out(and_512__out)
  );

  //Wire declarations for instance 'and_514' (Module coreir_and)
  wire [15:0] and_514__in0;
  wire [15:0] and_514__in1;
  wire [15:0] and_514__out;
  coreir_and #(.width(16)) and_514(
    .in0(and_514__in0),
    .in1(and_514__in1),
    .out(and_514__out)
  );

  //Wire declarations for instance 'and_516' (Module coreir_and)
  wire [15:0] and_516__in0;
  wire [15:0] and_516__in1;
  wire [15:0] and_516__out;
  coreir_and #(.width(16)) and_516(
    .in0(and_516__in0),
    .in1(and_516__in1),
    .out(and_516__out)
  );

  //Wire declarations for instance 'and_518' (Module coreir_and)
  wire [15:0] and_518__in0;
  wire [15:0] and_518__in1;
  wire [15:0] and_518__out;
  coreir_and #(.width(16)) and_518(
    .in0(and_518__in0),
    .in1(and_518__in1),
    .out(and_518__out)
  );

  //Wire declarations for instance 'and_52' (Module coreir_and)
  wire [15:0] and_52__in0;
  wire [15:0] and_52__in1;
  wire [15:0] and_52__out;
  coreir_and #(.width(16)) and_52(
    .in0(and_52__in0),
    .in1(and_52__in1),
    .out(and_52__out)
  );

  //Wire declarations for instance 'and_520' (Module coreir_and)
  wire [15:0] and_520__in0;
  wire [15:0] and_520__in1;
  wire [15:0] and_520__out;
  coreir_and #(.width(16)) and_520(
    .in0(and_520__in0),
    .in1(and_520__in1),
    .out(and_520__out)
  );

  //Wire declarations for instance 'and_522' (Module coreir_and)
  wire [15:0] and_522__in0;
  wire [15:0] and_522__in1;
  wire [15:0] and_522__out;
  coreir_and #(.width(16)) and_522(
    .in0(and_522__in0),
    .in1(and_522__in1),
    .out(and_522__out)
  );

  //Wire declarations for instance 'and_524' (Module coreir_and)
  wire [15:0] and_524__in0;
  wire [15:0] and_524__in1;
  wire [15:0] and_524__out;
  coreir_and #(.width(16)) and_524(
    .in0(and_524__in0),
    .in1(and_524__in1),
    .out(and_524__out)
  );

  //Wire declarations for instance 'and_526' (Module coreir_and)
  wire [15:0] and_526__in0;
  wire [15:0] and_526__in1;
  wire [15:0] and_526__out;
  coreir_and #(.width(16)) and_526(
    .in0(and_526__in0),
    .in1(and_526__in1),
    .out(and_526__out)
  );

  //Wire declarations for instance 'and_528' (Module coreir_and)
  wire [15:0] and_528__in0;
  wire [15:0] and_528__in1;
  wire [15:0] and_528__out;
  coreir_and #(.width(16)) and_528(
    .in0(and_528__in0),
    .in1(and_528__in1),
    .out(and_528__out)
  );

  //Wire declarations for instance 'and_530' (Module coreir_and)
  wire [15:0] and_530__in0;
  wire [15:0] and_530__in1;
  wire [15:0] and_530__out;
  coreir_and #(.width(16)) and_530(
    .in0(and_530__in0),
    .in1(and_530__in1),
    .out(and_530__out)
  );

  //Wire declarations for instance 'and_532' (Module coreir_and)
  wire [15:0] and_532__in0;
  wire [15:0] and_532__in1;
  wire [15:0] and_532__out;
  coreir_and #(.width(16)) and_532(
    .in0(and_532__in0),
    .in1(and_532__in1),
    .out(and_532__out)
  );

  //Wire declarations for instance 'and_534' (Module coreir_and)
  wire [15:0] and_534__in0;
  wire [15:0] and_534__in1;
  wire [15:0] and_534__out;
  coreir_and #(.width(16)) and_534(
    .in0(and_534__in0),
    .in1(and_534__in1),
    .out(and_534__out)
  );

  //Wire declarations for instance 'and_536' (Module coreir_and)
  wire [15:0] and_536__in0;
  wire [15:0] and_536__in1;
  wire [15:0] and_536__out;
  coreir_and #(.width(16)) and_536(
    .in0(and_536__in0),
    .in1(and_536__in1),
    .out(and_536__out)
  );

  //Wire declarations for instance 'and_538' (Module coreir_and)
  wire [15:0] and_538__in0;
  wire [15:0] and_538__in1;
  wire [15:0] and_538__out;
  coreir_and #(.width(16)) and_538(
    .in0(and_538__in0),
    .in1(and_538__in1),
    .out(and_538__out)
  );

  //Wire declarations for instance 'and_54' (Module coreir_and)
  wire [15:0] and_54__in0;
  wire [15:0] and_54__in1;
  wire [15:0] and_54__out;
  coreir_and #(.width(16)) and_54(
    .in0(and_54__in0),
    .in1(and_54__in1),
    .out(and_54__out)
  );

  //Wire declarations for instance 'and_540' (Module coreir_and)
  wire [15:0] and_540__in0;
  wire [15:0] and_540__in1;
  wire [15:0] and_540__out;
  coreir_and #(.width(16)) and_540(
    .in0(and_540__in0),
    .in1(and_540__in1),
    .out(and_540__out)
  );

  //Wire declarations for instance 'and_542' (Module coreir_and)
  wire [15:0] and_542__in0;
  wire [15:0] and_542__in1;
  wire [15:0] and_542__out;
  coreir_and #(.width(16)) and_542(
    .in0(and_542__in0),
    .in1(and_542__in1),
    .out(and_542__out)
  );

  //Wire declarations for instance 'and_544' (Module coreir_and)
  wire [15:0] and_544__in0;
  wire [15:0] and_544__in1;
  wire [15:0] and_544__out;
  coreir_and #(.width(16)) and_544(
    .in0(and_544__in0),
    .in1(and_544__in1),
    .out(and_544__out)
  );

  //Wire declarations for instance 'and_546' (Module coreir_and)
  wire [15:0] and_546__in0;
  wire [15:0] and_546__in1;
  wire [15:0] and_546__out;
  coreir_and #(.width(16)) and_546(
    .in0(and_546__in0),
    .in1(and_546__in1),
    .out(and_546__out)
  );

  //Wire declarations for instance 'and_548' (Module coreir_and)
  wire [15:0] and_548__in0;
  wire [15:0] and_548__in1;
  wire [15:0] and_548__out;
  coreir_and #(.width(16)) and_548(
    .in0(and_548__in0),
    .in1(and_548__in1),
    .out(and_548__out)
  );

  //Wire declarations for instance 'and_550' (Module coreir_and)
  wire [15:0] and_550__in0;
  wire [15:0] and_550__in1;
  wire [15:0] and_550__out;
  coreir_and #(.width(16)) and_550(
    .in0(and_550__in0),
    .in1(and_550__in1),
    .out(and_550__out)
  );

  //Wire declarations for instance 'and_552' (Module coreir_and)
  wire [15:0] and_552__in0;
  wire [15:0] and_552__in1;
  wire [15:0] and_552__out;
  coreir_and #(.width(16)) and_552(
    .in0(and_552__in0),
    .in1(and_552__in1),
    .out(and_552__out)
  );

  //Wire declarations for instance 'and_554' (Module coreir_and)
  wire [15:0] and_554__in0;
  wire [15:0] and_554__in1;
  wire [15:0] and_554__out;
  coreir_and #(.width(16)) and_554(
    .in0(and_554__in0),
    .in1(and_554__in1),
    .out(and_554__out)
  );

  //Wire declarations for instance 'and_556' (Module coreir_and)
  wire [15:0] and_556__in0;
  wire [15:0] and_556__in1;
  wire [15:0] and_556__out;
  coreir_and #(.width(16)) and_556(
    .in0(and_556__in0),
    .in1(and_556__in1),
    .out(and_556__out)
  );

  //Wire declarations for instance 'and_558' (Module coreir_and)
  wire [15:0] and_558__in0;
  wire [15:0] and_558__in1;
  wire [15:0] and_558__out;
  coreir_and #(.width(16)) and_558(
    .in0(and_558__in0),
    .in1(and_558__in1),
    .out(and_558__out)
  );

  //Wire declarations for instance 'and_56' (Module coreir_and)
  wire [15:0] and_56__in0;
  wire [15:0] and_56__in1;
  wire [15:0] and_56__out;
  coreir_and #(.width(16)) and_56(
    .in0(and_56__in0),
    .in1(and_56__in1),
    .out(and_56__out)
  );

  //Wire declarations for instance 'and_560' (Module coreir_and)
  wire [15:0] and_560__in0;
  wire [15:0] and_560__in1;
  wire [15:0] and_560__out;
  coreir_and #(.width(16)) and_560(
    .in0(and_560__in0),
    .in1(and_560__in1),
    .out(and_560__out)
  );

  //Wire declarations for instance 'and_562' (Module coreir_and)
  wire [15:0] and_562__in0;
  wire [15:0] and_562__in1;
  wire [15:0] and_562__out;
  coreir_and #(.width(16)) and_562(
    .in0(and_562__in0),
    .in1(and_562__in1),
    .out(and_562__out)
  );

  //Wire declarations for instance 'and_564' (Module coreir_and)
  wire [15:0] and_564__in0;
  wire [15:0] and_564__in1;
  wire [15:0] and_564__out;
  coreir_and #(.width(16)) and_564(
    .in0(and_564__in0),
    .in1(and_564__in1),
    .out(and_564__out)
  );

  //Wire declarations for instance 'and_566' (Module coreir_and)
  wire [15:0] and_566__in0;
  wire [15:0] and_566__in1;
  wire [15:0] and_566__out;
  coreir_and #(.width(16)) and_566(
    .in0(and_566__in0),
    .in1(and_566__in1),
    .out(and_566__out)
  );

  //Wire declarations for instance 'and_568' (Module coreir_and)
  wire [15:0] and_568__in0;
  wire [15:0] and_568__in1;
  wire [15:0] and_568__out;
  coreir_and #(.width(16)) and_568(
    .in0(and_568__in0),
    .in1(and_568__in1),
    .out(and_568__out)
  );

  //Wire declarations for instance 'and_570' (Module coreir_and)
  wire [15:0] and_570__in0;
  wire [15:0] and_570__in1;
  wire [15:0] and_570__out;
  coreir_and #(.width(16)) and_570(
    .in0(and_570__in0),
    .in1(and_570__in1),
    .out(and_570__out)
  );

  //Wire declarations for instance 'and_572' (Module coreir_and)
  wire [15:0] and_572__in0;
  wire [15:0] and_572__in1;
  wire [15:0] and_572__out;
  coreir_and #(.width(16)) and_572(
    .in0(and_572__in0),
    .in1(and_572__in1),
    .out(and_572__out)
  );

  //Wire declarations for instance 'and_574' (Module coreir_and)
  wire [15:0] and_574__in0;
  wire [15:0] and_574__in1;
  wire [15:0] and_574__out;
  coreir_and #(.width(16)) and_574(
    .in0(and_574__in0),
    .in1(and_574__in1),
    .out(and_574__out)
  );

  //Wire declarations for instance 'and_576' (Module coreir_and)
  wire [15:0] and_576__in0;
  wire [15:0] and_576__in1;
  wire [15:0] and_576__out;
  coreir_and #(.width(16)) and_576(
    .in0(and_576__in0),
    .in1(and_576__in1),
    .out(and_576__out)
  );

  //Wire declarations for instance 'and_578' (Module coreir_and)
  wire [15:0] and_578__in0;
  wire [15:0] and_578__in1;
  wire [15:0] and_578__out;
  coreir_and #(.width(16)) and_578(
    .in0(and_578__in0),
    .in1(and_578__in1),
    .out(and_578__out)
  );

  //Wire declarations for instance 'and_58' (Module coreir_and)
  wire [15:0] and_58__in0;
  wire [15:0] and_58__in1;
  wire [15:0] and_58__out;
  coreir_and #(.width(16)) and_58(
    .in0(and_58__in0),
    .in1(and_58__in1),
    .out(and_58__out)
  );

  //Wire declarations for instance 'and_580' (Module coreir_and)
  wire [15:0] and_580__in0;
  wire [15:0] and_580__in1;
  wire [15:0] and_580__out;
  coreir_and #(.width(16)) and_580(
    .in0(and_580__in0),
    .in1(and_580__in1),
    .out(and_580__out)
  );

  //Wire declarations for instance 'and_582' (Module coreir_and)
  wire [15:0] and_582__in0;
  wire [15:0] and_582__in1;
  wire [15:0] and_582__out;
  coreir_and #(.width(16)) and_582(
    .in0(and_582__in0),
    .in1(and_582__in1),
    .out(and_582__out)
  );

  //Wire declarations for instance 'and_584' (Module coreir_and)
  wire [15:0] and_584__in0;
  wire [15:0] and_584__in1;
  wire [15:0] and_584__out;
  coreir_and #(.width(16)) and_584(
    .in0(and_584__in0),
    .in1(and_584__in1),
    .out(and_584__out)
  );

  //Wire declarations for instance 'and_586' (Module coreir_and)
  wire [15:0] and_586__in0;
  wire [15:0] and_586__in1;
  wire [15:0] and_586__out;
  coreir_and #(.width(16)) and_586(
    .in0(and_586__in0),
    .in1(and_586__in1),
    .out(and_586__out)
  );

  //Wire declarations for instance 'and_588' (Module coreir_and)
  wire [15:0] and_588__in0;
  wire [15:0] and_588__in1;
  wire [15:0] and_588__out;
  coreir_and #(.width(16)) and_588(
    .in0(and_588__in0),
    .in1(and_588__in1),
    .out(and_588__out)
  );

  //Wire declarations for instance 'and_590' (Module coreir_and)
  wire [15:0] and_590__in0;
  wire [15:0] and_590__in1;
  wire [15:0] and_590__out;
  coreir_and #(.width(16)) and_590(
    .in0(and_590__in0),
    .in1(and_590__in1),
    .out(and_590__out)
  );

  //Wire declarations for instance 'and_592' (Module coreir_and)
  wire [15:0] and_592__in0;
  wire [15:0] and_592__in1;
  wire [15:0] and_592__out;
  coreir_and #(.width(16)) and_592(
    .in0(and_592__in0),
    .in1(and_592__in1),
    .out(and_592__out)
  );

  //Wire declarations for instance 'and_594' (Module coreir_and)
  wire [15:0] and_594__in0;
  wire [15:0] and_594__in1;
  wire [15:0] and_594__out;
  coreir_and #(.width(16)) and_594(
    .in0(and_594__in0),
    .in1(and_594__in1),
    .out(and_594__out)
  );

  //Wire declarations for instance 'and_596' (Module coreir_and)
  wire [15:0] and_596__in0;
  wire [15:0] and_596__in1;
  wire [15:0] and_596__out;
  coreir_and #(.width(16)) and_596(
    .in0(and_596__in0),
    .in1(and_596__in1),
    .out(and_596__out)
  );

  //Wire declarations for instance 'and_598' (Module coreir_and)
  wire [15:0] and_598__in0;
  wire [15:0] and_598__in1;
  wire [15:0] and_598__out;
  coreir_and #(.width(16)) and_598(
    .in0(and_598__in0),
    .in1(and_598__in1),
    .out(and_598__out)
  );

  //Wire declarations for instance 'and_6' (Module coreir_and)
  wire [15:0] and_6__in0;
  wire [15:0] and_6__in1;
  wire [15:0] and_6__out;
  coreir_and #(.width(16)) and_6(
    .in0(and_6__in0),
    .in1(and_6__in1),
    .out(and_6__out)
  );

  //Wire declarations for instance 'and_60' (Module coreir_and)
  wire [15:0] and_60__in0;
  wire [15:0] and_60__in1;
  wire [15:0] and_60__out;
  coreir_and #(.width(16)) and_60(
    .in0(and_60__in0),
    .in1(and_60__in1),
    .out(and_60__out)
  );

  //Wire declarations for instance 'and_600' (Module coreir_and)
  wire [15:0] and_600__in0;
  wire [15:0] and_600__in1;
  wire [15:0] and_600__out;
  coreir_and #(.width(16)) and_600(
    .in0(and_600__in0),
    .in1(and_600__in1),
    .out(and_600__out)
  );

  //Wire declarations for instance 'and_602' (Module coreir_and)
  wire [15:0] and_602__in0;
  wire [15:0] and_602__in1;
  wire [15:0] and_602__out;
  coreir_and #(.width(16)) and_602(
    .in0(and_602__in0),
    .in1(and_602__in1),
    .out(and_602__out)
  );

  //Wire declarations for instance 'and_604' (Module coreir_and)
  wire [15:0] and_604__in0;
  wire [15:0] and_604__in1;
  wire [15:0] and_604__out;
  coreir_and #(.width(16)) and_604(
    .in0(and_604__in0),
    .in1(and_604__in1),
    .out(and_604__out)
  );

  //Wire declarations for instance 'and_606' (Module coreir_and)
  wire [15:0] and_606__in0;
  wire [15:0] and_606__in1;
  wire [15:0] and_606__out;
  coreir_and #(.width(16)) and_606(
    .in0(and_606__in0),
    .in1(and_606__in1),
    .out(and_606__out)
  );

  //Wire declarations for instance 'and_608' (Module coreir_and)
  wire [15:0] and_608__in0;
  wire [15:0] and_608__in1;
  wire [15:0] and_608__out;
  coreir_and #(.width(16)) and_608(
    .in0(and_608__in0),
    .in1(and_608__in1),
    .out(and_608__out)
  );

  //Wire declarations for instance 'and_610' (Module coreir_and)
  wire [15:0] and_610__in0;
  wire [15:0] and_610__in1;
  wire [15:0] and_610__out;
  coreir_and #(.width(16)) and_610(
    .in0(and_610__in0),
    .in1(and_610__in1),
    .out(and_610__out)
  );

  //Wire declarations for instance 'and_612' (Module coreir_and)
  wire [15:0] and_612__in0;
  wire [15:0] and_612__in1;
  wire [15:0] and_612__out;
  coreir_and #(.width(16)) and_612(
    .in0(and_612__in0),
    .in1(and_612__in1),
    .out(and_612__out)
  );

  //Wire declarations for instance 'and_614' (Module coreir_and)
  wire [15:0] and_614__in0;
  wire [15:0] and_614__in1;
  wire [15:0] and_614__out;
  coreir_and #(.width(16)) and_614(
    .in0(and_614__in0),
    .in1(and_614__in1),
    .out(and_614__out)
  );

  //Wire declarations for instance 'and_616' (Module coreir_and)
  wire [15:0] and_616__in0;
  wire [15:0] and_616__in1;
  wire [15:0] and_616__out;
  coreir_and #(.width(16)) and_616(
    .in0(and_616__in0),
    .in1(and_616__in1),
    .out(and_616__out)
  );

  //Wire declarations for instance 'and_618' (Module coreir_and)
  wire [15:0] and_618__in0;
  wire [15:0] and_618__in1;
  wire [15:0] and_618__out;
  coreir_and #(.width(16)) and_618(
    .in0(and_618__in0),
    .in1(and_618__in1),
    .out(and_618__out)
  );

  //Wire declarations for instance 'and_62' (Module coreir_and)
  wire [15:0] and_62__in0;
  wire [15:0] and_62__in1;
  wire [15:0] and_62__out;
  coreir_and #(.width(16)) and_62(
    .in0(and_62__in0),
    .in1(and_62__in1),
    .out(and_62__out)
  );

  //Wire declarations for instance 'and_620' (Module coreir_and)
  wire [15:0] and_620__in0;
  wire [15:0] and_620__in1;
  wire [15:0] and_620__out;
  coreir_and #(.width(16)) and_620(
    .in0(and_620__in0),
    .in1(and_620__in1),
    .out(and_620__out)
  );

  //Wire declarations for instance 'and_622' (Module coreir_and)
  wire [15:0] and_622__in0;
  wire [15:0] and_622__in1;
  wire [15:0] and_622__out;
  coreir_and #(.width(16)) and_622(
    .in0(and_622__in0),
    .in1(and_622__in1),
    .out(and_622__out)
  );

  //Wire declarations for instance 'and_624' (Module coreir_and)
  wire [15:0] and_624__in0;
  wire [15:0] and_624__in1;
  wire [15:0] and_624__out;
  coreir_and #(.width(16)) and_624(
    .in0(and_624__in0),
    .in1(and_624__in1),
    .out(and_624__out)
  );

  //Wire declarations for instance 'and_626' (Module coreir_and)
  wire [15:0] and_626__in0;
  wire [15:0] and_626__in1;
  wire [15:0] and_626__out;
  coreir_and #(.width(16)) and_626(
    .in0(and_626__in0),
    .in1(and_626__in1),
    .out(and_626__out)
  );

  //Wire declarations for instance 'and_628' (Module coreir_and)
  wire [15:0] and_628__in0;
  wire [15:0] and_628__in1;
  wire [15:0] and_628__out;
  coreir_and #(.width(16)) and_628(
    .in0(and_628__in0),
    .in1(and_628__in1),
    .out(and_628__out)
  );

  //Wire declarations for instance 'and_630' (Module coreir_and)
  wire [15:0] and_630__in0;
  wire [15:0] and_630__in1;
  wire [15:0] and_630__out;
  coreir_and #(.width(16)) and_630(
    .in0(and_630__in0),
    .in1(and_630__in1),
    .out(and_630__out)
  );

  //Wire declarations for instance 'and_632' (Module coreir_and)
  wire [15:0] and_632__in0;
  wire [15:0] and_632__in1;
  wire [15:0] and_632__out;
  coreir_and #(.width(16)) and_632(
    .in0(and_632__in0),
    .in1(and_632__in1),
    .out(and_632__out)
  );

  //Wire declarations for instance 'and_634' (Module coreir_and)
  wire [15:0] and_634__in0;
  wire [15:0] and_634__in1;
  wire [15:0] and_634__out;
  coreir_and #(.width(16)) and_634(
    .in0(and_634__in0),
    .in1(and_634__in1),
    .out(and_634__out)
  );

  //Wire declarations for instance 'and_636' (Module coreir_and)
  wire [15:0] and_636__in0;
  wire [15:0] and_636__in1;
  wire [15:0] and_636__out;
  coreir_and #(.width(16)) and_636(
    .in0(and_636__in0),
    .in1(and_636__in1),
    .out(and_636__out)
  );

  //Wire declarations for instance 'and_638' (Module coreir_and)
  wire [15:0] and_638__in0;
  wire [15:0] and_638__in1;
  wire [15:0] and_638__out;
  coreir_and #(.width(16)) and_638(
    .in0(and_638__in0),
    .in1(and_638__in1),
    .out(and_638__out)
  );

  //Wire declarations for instance 'and_64' (Module coreir_and)
  wire [15:0] and_64__in0;
  wire [15:0] and_64__in1;
  wire [15:0] and_64__out;
  coreir_and #(.width(16)) and_64(
    .in0(and_64__in0),
    .in1(and_64__in1),
    .out(and_64__out)
  );

  //Wire declarations for instance 'and_640' (Module coreir_and)
  wire [15:0] and_640__in0;
  wire [15:0] and_640__in1;
  wire [15:0] and_640__out;
  coreir_and #(.width(16)) and_640(
    .in0(and_640__in0),
    .in1(and_640__in1),
    .out(and_640__out)
  );

  //Wire declarations for instance 'and_642' (Module coreir_and)
  wire [15:0] and_642__in0;
  wire [15:0] and_642__in1;
  wire [15:0] and_642__out;
  coreir_and #(.width(16)) and_642(
    .in0(and_642__in0),
    .in1(and_642__in1),
    .out(and_642__out)
  );

  //Wire declarations for instance 'and_644' (Module coreir_and)
  wire [15:0] and_644__in0;
  wire [15:0] and_644__in1;
  wire [15:0] and_644__out;
  coreir_and #(.width(16)) and_644(
    .in0(and_644__in0),
    .in1(and_644__in1),
    .out(and_644__out)
  );

  //Wire declarations for instance 'and_646' (Module coreir_and)
  wire [15:0] and_646__in0;
  wire [15:0] and_646__in1;
  wire [15:0] and_646__out;
  coreir_and #(.width(16)) and_646(
    .in0(and_646__in0),
    .in1(and_646__in1),
    .out(and_646__out)
  );

  //Wire declarations for instance 'and_648' (Module coreir_and)
  wire [15:0] and_648__in0;
  wire [15:0] and_648__in1;
  wire [15:0] and_648__out;
  coreir_and #(.width(16)) and_648(
    .in0(and_648__in0),
    .in1(and_648__in1),
    .out(and_648__out)
  );

  //Wire declarations for instance 'and_650' (Module coreir_and)
  wire [15:0] and_650__in0;
  wire [15:0] and_650__in1;
  wire [15:0] and_650__out;
  coreir_and #(.width(16)) and_650(
    .in0(and_650__in0),
    .in1(and_650__in1),
    .out(and_650__out)
  );

  //Wire declarations for instance 'and_652' (Module coreir_and)
  wire [15:0] and_652__in0;
  wire [15:0] and_652__in1;
  wire [15:0] and_652__out;
  coreir_and #(.width(16)) and_652(
    .in0(and_652__in0),
    .in1(and_652__in1),
    .out(and_652__out)
  );

  //Wire declarations for instance 'and_654' (Module coreir_and)
  wire [15:0] and_654__in0;
  wire [15:0] and_654__in1;
  wire [15:0] and_654__out;
  coreir_and #(.width(16)) and_654(
    .in0(and_654__in0),
    .in1(and_654__in1),
    .out(and_654__out)
  );

  //Wire declarations for instance 'and_656' (Module coreir_and)
  wire [15:0] and_656__in0;
  wire [15:0] and_656__in1;
  wire [15:0] and_656__out;
  coreir_and #(.width(16)) and_656(
    .in0(and_656__in0),
    .in1(and_656__in1),
    .out(and_656__out)
  );

  //Wire declarations for instance 'and_658' (Module coreir_and)
  wire [15:0] and_658__in0;
  wire [15:0] and_658__in1;
  wire [15:0] and_658__out;
  coreir_and #(.width(16)) and_658(
    .in0(and_658__in0),
    .in1(and_658__in1),
    .out(and_658__out)
  );

  //Wire declarations for instance 'and_66' (Module coreir_and)
  wire [15:0] and_66__in0;
  wire [15:0] and_66__in1;
  wire [15:0] and_66__out;
  coreir_and #(.width(16)) and_66(
    .in0(and_66__in0),
    .in1(and_66__in1),
    .out(and_66__out)
  );

  //Wire declarations for instance 'and_660' (Module coreir_and)
  wire [15:0] and_660__in0;
  wire [15:0] and_660__in1;
  wire [15:0] and_660__out;
  coreir_and #(.width(16)) and_660(
    .in0(and_660__in0),
    .in1(and_660__in1),
    .out(and_660__out)
  );

  //Wire declarations for instance 'and_662' (Module coreir_and)
  wire [15:0] and_662__in0;
  wire [15:0] and_662__in1;
  wire [15:0] and_662__out;
  coreir_and #(.width(16)) and_662(
    .in0(and_662__in0),
    .in1(and_662__in1),
    .out(and_662__out)
  );

  //Wire declarations for instance 'and_664' (Module coreir_and)
  wire [15:0] and_664__in0;
  wire [15:0] and_664__in1;
  wire [15:0] and_664__out;
  coreir_and #(.width(16)) and_664(
    .in0(and_664__in0),
    .in1(and_664__in1),
    .out(and_664__out)
  );

  //Wire declarations for instance 'and_666' (Module coreir_and)
  wire [15:0] and_666__in0;
  wire [15:0] and_666__in1;
  wire [15:0] and_666__out;
  coreir_and #(.width(16)) and_666(
    .in0(and_666__in0),
    .in1(and_666__in1),
    .out(and_666__out)
  );

  //Wire declarations for instance 'and_668' (Module coreir_and)
  wire [15:0] and_668__in0;
  wire [15:0] and_668__in1;
  wire [15:0] and_668__out;
  coreir_and #(.width(16)) and_668(
    .in0(and_668__in0),
    .in1(and_668__in1),
    .out(and_668__out)
  );

  //Wire declarations for instance 'and_670' (Module coreir_and)
  wire [15:0] and_670__in0;
  wire [15:0] and_670__in1;
  wire [15:0] and_670__out;
  coreir_and #(.width(16)) and_670(
    .in0(and_670__in0),
    .in1(and_670__in1),
    .out(and_670__out)
  );

  //Wire declarations for instance 'and_672' (Module coreir_and)
  wire [15:0] and_672__in0;
  wire [15:0] and_672__in1;
  wire [15:0] and_672__out;
  coreir_and #(.width(16)) and_672(
    .in0(and_672__in0),
    .in1(and_672__in1),
    .out(and_672__out)
  );

  //Wire declarations for instance 'and_674' (Module coreir_and)
  wire [15:0] and_674__in0;
  wire [15:0] and_674__in1;
  wire [15:0] and_674__out;
  coreir_and #(.width(16)) and_674(
    .in0(and_674__in0),
    .in1(and_674__in1),
    .out(and_674__out)
  );

  //Wire declarations for instance 'and_676' (Module coreir_and)
  wire [15:0] and_676__in0;
  wire [15:0] and_676__in1;
  wire [15:0] and_676__out;
  coreir_and #(.width(16)) and_676(
    .in0(and_676__in0),
    .in1(and_676__in1),
    .out(and_676__out)
  );

  //Wire declarations for instance 'and_678' (Module coreir_and)
  wire [15:0] and_678__in0;
  wire [15:0] and_678__in1;
  wire [15:0] and_678__out;
  coreir_and #(.width(16)) and_678(
    .in0(and_678__in0),
    .in1(and_678__in1),
    .out(and_678__out)
  );

  //Wire declarations for instance 'and_68' (Module coreir_and)
  wire [15:0] and_68__in0;
  wire [15:0] and_68__in1;
  wire [15:0] and_68__out;
  coreir_and #(.width(16)) and_68(
    .in0(and_68__in0),
    .in1(and_68__in1),
    .out(and_68__out)
  );

  //Wire declarations for instance 'and_680' (Module coreir_and)
  wire [15:0] and_680__in0;
  wire [15:0] and_680__in1;
  wire [15:0] and_680__out;
  coreir_and #(.width(16)) and_680(
    .in0(and_680__in0),
    .in1(and_680__in1),
    .out(and_680__out)
  );

  //Wire declarations for instance 'and_682' (Module coreir_and)
  wire [15:0] and_682__in0;
  wire [15:0] and_682__in1;
  wire [15:0] and_682__out;
  coreir_and #(.width(16)) and_682(
    .in0(and_682__in0),
    .in1(and_682__in1),
    .out(and_682__out)
  );

  //Wire declarations for instance 'and_684' (Module coreir_and)
  wire [15:0] and_684__in0;
  wire [15:0] and_684__in1;
  wire [15:0] and_684__out;
  coreir_and #(.width(16)) and_684(
    .in0(and_684__in0),
    .in1(and_684__in1),
    .out(and_684__out)
  );

  //Wire declarations for instance 'and_686' (Module coreir_and)
  wire [15:0] and_686__in0;
  wire [15:0] and_686__in1;
  wire [15:0] and_686__out;
  coreir_and #(.width(16)) and_686(
    .in0(and_686__in0),
    .in1(and_686__in1),
    .out(and_686__out)
  );

  //Wire declarations for instance 'and_688' (Module coreir_and)
  wire [15:0] and_688__in0;
  wire [15:0] and_688__in1;
  wire [15:0] and_688__out;
  coreir_and #(.width(16)) and_688(
    .in0(and_688__in0),
    .in1(and_688__in1),
    .out(and_688__out)
  );

  //Wire declarations for instance 'and_690' (Module coreir_and)
  wire [15:0] and_690__in0;
  wire [15:0] and_690__in1;
  wire [15:0] and_690__out;
  coreir_and #(.width(16)) and_690(
    .in0(and_690__in0),
    .in1(and_690__in1),
    .out(and_690__out)
  );

  //Wire declarations for instance 'and_692' (Module coreir_and)
  wire [15:0] and_692__in0;
  wire [15:0] and_692__in1;
  wire [15:0] and_692__out;
  coreir_and #(.width(16)) and_692(
    .in0(and_692__in0),
    .in1(and_692__in1),
    .out(and_692__out)
  );

  //Wire declarations for instance 'and_694' (Module coreir_and)
  wire [15:0] and_694__in0;
  wire [15:0] and_694__in1;
  wire [15:0] and_694__out;
  coreir_and #(.width(16)) and_694(
    .in0(and_694__in0),
    .in1(and_694__in1),
    .out(and_694__out)
  );

  //Wire declarations for instance 'and_696' (Module coreir_and)
  wire [15:0] and_696__in0;
  wire [15:0] and_696__in1;
  wire [15:0] and_696__out;
  coreir_and #(.width(16)) and_696(
    .in0(and_696__in0),
    .in1(and_696__in1),
    .out(and_696__out)
  );

  //Wire declarations for instance 'and_698' (Module coreir_and)
  wire [15:0] and_698__in0;
  wire [15:0] and_698__in1;
  wire [15:0] and_698__out;
  coreir_and #(.width(16)) and_698(
    .in0(and_698__in0),
    .in1(and_698__in1),
    .out(and_698__out)
  );

  //Wire declarations for instance 'and_70' (Module coreir_and)
  wire [15:0] and_70__in0;
  wire [15:0] and_70__in1;
  wire [15:0] and_70__out;
  coreir_and #(.width(16)) and_70(
    .in0(and_70__in0),
    .in1(and_70__in1),
    .out(and_70__out)
  );

  //Wire declarations for instance 'and_700' (Module coreir_and)
  wire [15:0] and_700__in0;
  wire [15:0] and_700__in1;
  wire [15:0] and_700__out;
  coreir_and #(.width(16)) and_700(
    .in0(and_700__in0),
    .in1(and_700__in1),
    .out(and_700__out)
  );

  //Wire declarations for instance 'and_702' (Module coreir_and)
  wire [15:0] and_702__in0;
  wire [15:0] and_702__in1;
  wire [15:0] and_702__out;
  coreir_and #(.width(16)) and_702(
    .in0(and_702__in0),
    .in1(and_702__in1),
    .out(and_702__out)
  );

  //Wire declarations for instance 'and_704' (Module coreir_and)
  wire [15:0] and_704__in0;
  wire [15:0] and_704__in1;
  wire [15:0] and_704__out;
  coreir_and #(.width(16)) and_704(
    .in0(and_704__in0),
    .in1(and_704__in1),
    .out(and_704__out)
  );

  //Wire declarations for instance 'and_706' (Module coreir_and)
  wire [15:0] and_706__in0;
  wire [15:0] and_706__in1;
  wire [15:0] and_706__out;
  coreir_and #(.width(16)) and_706(
    .in0(and_706__in0),
    .in1(and_706__in1),
    .out(and_706__out)
  );

  //Wire declarations for instance 'and_708' (Module coreir_and)
  wire [15:0] and_708__in0;
  wire [15:0] and_708__in1;
  wire [15:0] and_708__out;
  coreir_and #(.width(16)) and_708(
    .in0(and_708__in0),
    .in1(and_708__in1),
    .out(and_708__out)
  );

  //Wire declarations for instance 'and_710' (Module coreir_and)
  wire [15:0] and_710__in0;
  wire [15:0] and_710__in1;
  wire [15:0] and_710__out;
  coreir_and #(.width(16)) and_710(
    .in0(and_710__in0),
    .in1(and_710__in1),
    .out(and_710__out)
  );

  //Wire declarations for instance 'and_712' (Module coreir_and)
  wire [15:0] and_712__in0;
  wire [15:0] and_712__in1;
  wire [15:0] and_712__out;
  coreir_and #(.width(16)) and_712(
    .in0(and_712__in0),
    .in1(and_712__in1),
    .out(and_712__out)
  );

  //Wire declarations for instance 'and_714' (Module coreir_and)
  wire [15:0] and_714__in0;
  wire [15:0] and_714__in1;
  wire [15:0] and_714__out;
  coreir_and #(.width(16)) and_714(
    .in0(and_714__in0),
    .in1(and_714__in1),
    .out(and_714__out)
  );

  //Wire declarations for instance 'and_716' (Module coreir_and)
  wire [15:0] and_716__in0;
  wire [15:0] and_716__in1;
  wire [15:0] and_716__out;
  coreir_and #(.width(16)) and_716(
    .in0(and_716__in0),
    .in1(and_716__in1),
    .out(and_716__out)
  );

  //Wire declarations for instance 'and_718' (Module coreir_and)
  wire [15:0] and_718__in0;
  wire [15:0] and_718__in1;
  wire [15:0] and_718__out;
  coreir_and #(.width(16)) and_718(
    .in0(and_718__in0),
    .in1(and_718__in1),
    .out(and_718__out)
  );

  //Wire declarations for instance 'and_72' (Module coreir_and)
  wire [15:0] and_72__in0;
  wire [15:0] and_72__in1;
  wire [15:0] and_72__out;
  coreir_and #(.width(16)) and_72(
    .in0(and_72__in0),
    .in1(and_72__in1),
    .out(and_72__out)
  );

  //Wire declarations for instance 'and_720' (Module coreir_and)
  wire [15:0] and_720__in0;
  wire [15:0] and_720__in1;
  wire [15:0] and_720__out;
  coreir_and #(.width(16)) and_720(
    .in0(and_720__in0),
    .in1(and_720__in1),
    .out(and_720__out)
  );

  //Wire declarations for instance 'and_722' (Module coreir_and)
  wire [15:0] and_722__in0;
  wire [15:0] and_722__in1;
  wire [15:0] and_722__out;
  coreir_and #(.width(16)) and_722(
    .in0(and_722__in0),
    .in1(and_722__in1),
    .out(and_722__out)
  );

  //Wire declarations for instance 'and_724' (Module coreir_and)
  wire [15:0] and_724__in0;
  wire [15:0] and_724__in1;
  wire [15:0] and_724__out;
  coreir_and #(.width(16)) and_724(
    .in0(and_724__in0),
    .in1(and_724__in1),
    .out(and_724__out)
  );

  //Wire declarations for instance 'and_726' (Module coreir_and)
  wire [15:0] and_726__in0;
  wire [15:0] and_726__in1;
  wire [15:0] and_726__out;
  coreir_and #(.width(16)) and_726(
    .in0(and_726__in0),
    .in1(and_726__in1),
    .out(and_726__out)
  );

  //Wire declarations for instance 'and_728' (Module coreir_and)
  wire [15:0] and_728__in0;
  wire [15:0] and_728__in1;
  wire [15:0] and_728__out;
  coreir_and #(.width(16)) and_728(
    .in0(and_728__in0),
    .in1(and_728__in1),
    .out(and_728__out)
  );

  //Wire declarations for instance 'and_730' (Module coreir_and)
  wire [15:0] and_730__in0;
  wire [15:0] and_730__in1;
  wire [15:0] and_730__out;
  coreir_and #(.width(16)) and_730(
    .in0(and_730__in0),
    .in1(and_730__in1),
    .out(and_730__out)
  );

  //Wire declarations for instance 'and_732' (Module coreir_and)
  wire [15:0] and_732__in0;
  wire [15:0] and_732__in1;
  wire [15:0] and_732__out;
  coreir_and #(.width(16)) and_732(
    .in0(and_732__in0),
    .in1(and_732__in1),
    .out(and_732__out)
  );

  //Wire declarations for instance 'and_734' (Module coreir_and)
  wire [15:0] and_734__in0;
  wire [15:0] and_734__in1;
  wire [15:0] and_734__out;
  coreir_and #(.width(16)) and_734(
    .in0(and_734__in0),
    .in1(and_734__in1),
    .out(and_734__out)
  );

  //Wire declarations for instance 'and_736' (Module coreir_and)
  wire [15:0] and_736__in0;
  wire [15:0] and_736__in1;
  wire [15:0] and_736__out;
  coreir_and #(.width(16)) and_736(
    .in0(and_736__in0),
    .in1(and_736__in1),
    .out(and_736__out)
  );

  //Wire declarations for instance 'and_738' (Module coreir_and)
  wire [15:0] and_738__in0;
  wire [15:0] and_738__in1;
  wire [15:0] and_738__out;
  coreir_and #(.width(16)) and_738(
    .in0(and_738__in0),
    .in1(and_738__in1),
    .out(and_738__out)
  );

  //Wire declarations for instance 'and_74' (Module coreir_and)
  wire [15:0] and_74__in0;
  wire [15:0] and_74__in1;
  wire [15:0] and_74__out;
  coreir_and #(.width(16)) and_74(
    .in0(and_74__in0),
    .in1(and_74__in1),
    .out(and_74__out)
  );

  //Wire declarations for instance 'and_740' (Module coreir_and)
  wire [15:0] and_740__in0;
  wire [15:0] and_740__in1;
  wire [15:0] and_740__out;
  coreir_and #(.width(16)) and_740(
    .in0(and_740__in0),
    .in1(and_740__in1),
    .out(and_740__out)
  );

  //Wire declarations for instance 'and_742' (Module coreir_and)
  wire [15:0] and_742__in0;
  wire [15:0] and_742__in1;
  wire [15:0] and_742__out;
  coreir_and #(.width(16)) and_742(
    .in0(and_742__in0),
    .in1(and_742__in1),
    .out(and_742__out)
  );

  //Wire declarations for instance 'and_744' (Module coreir_and)
  wire [15:0] and_744__in0;
  wire [15:0] and_744__in1;
  wire [15:0] and_744__out;
  coreir_and #(.width(16)) and_744(
    .in0(and_744__in0),
    .in1(and_744__in1),
    .out(and_744__out)
  );

  //Wire declarations for instance 'and_746' (Module coreir_and)
  wire [15:0] and_746__in0;
  wire [15:0] and_746__in1;
  wire [15:0] and_746__out;
  coreir_and #(.width(16)) and_746(
    .in0(and_746__in0),
    .in1(and_746__in1),
    .out(and_746__out)
  );

  //Wire declarations for instance 'and_748' (Module coreir_and)
  wire [15:0] and_748__in0;
  wire [15:0] and_748__in1;
  wire [15:0] and_748__out;
  coreir_and #(.width(16)) and_748(
    .in0(and_748__in0),
    .in1(and_748__in1),
    .out(and_748__out)
  );

  //Wire declarations for instance 'and_750' (Module coreir_and)
  wire [15:0] and_750__in0;
  wire [15:0] and_750__in1;
  wire [15:0] and_750__out;
  coreir_and #(.width(16)) and_750(
    .in0(and_750__in0),
    .in1(and_750__in1),
    .out(and_750__out)
  );

  //Wire declarations for instance 'and_752' (Module coreir_and)
  wire [15:0] and_752__in0;
  wire [15:0] and_752__in1;
  wire [15:0] and_752__out;
  coreir_and #(.width(16)) and_752(
    .in0(and_752__in0),
    .in1(and_752__in1),
    .out(and_752__out)
  );

  //Wire declarations for instance 'and_754' (Module coreir_and)
  wire [15:0] and_754__in0;
  wire [15:0] and_754__in1;
  wire [15:0] and_754__out;
  coreir_and #(.width(16)) and_754(
    .in0(and_754__in0),
    .in1(and_754__in1),
    .out(and_754__out)
  );

  //Wire declarations for instance 'and_756' (Module coreir_and)
  wire [15:0] and_756__in0;
  wire [15:0] and_756__in1;
  wire [15:0] and_756__out;
  coreir_and #(.width(16)) and_756(
    .in0(and_756__in0),
    .in1(and_756__in1),
    .out(and_756__out)
  );

  //Wire declarations for instance 'and_758' (Module coreir_and)
  wire [15:0] and_758__in0;
  wire [15:0] and_758__in1;
  wire [15:0] and_758__out;
  coreir_and #(.width(16)) and_758(
    .in0(and_758__in0),
    .in1(and_758__in1),
    .out(and_758__out)
  );

  //Wire declarations for instance 'and_76' (Module coreir_and)
  wire [15:0] and_76__in0;
  wire [15:0] and_76__in1;
  wire [15:0] and_76__out;
  coreir_and #(.width(16)) and_76(
    .in0(and_76__in0),
    .in1(and_76__in1),
    .out(and_76__out)
  );

  //Wire declarations for instance 'and_760' (Module coreir_and)
  wire [15:0] and_760__in0;
  wire [15:0] and_760__in1;
  wire [15:0] and_760__out;
  coreir_and #(.width(16)) and_760(
    .in0(and_760__in0),
    .in1(and_760__in1),
    .out(and_760__out)
  );

  //Wire declarations for instance 'and_762' (Module coreir_and)
  wire [15:0] and_762__in0;
  wire [15:0] and_762__in1;
  wire [15:0] and_762__out;
  coreir_and #(.width(16)) and_762(
    .in0(and_762__in0),
    .in1(and_762__in1),
    .out(and_762__out)
  );

  //Wire declarations for instance 'and_764' (Module coreir_and)
  wire [15:0] and_764__in0;
  wire [15:0] and_764__in1;
  wire [15:0] and_764__out;
  coreir_and #(.width(16)) and_764(
    .in0(and_764__in0),
    .in1(and_764__in1),
    .out(and_764__out)
  );

  //Wire declarations for instance 'and_766' (Module coreir_and)
  wire [15:0] and_766__in0;
  wire [15:0] and_766__in1;
  wire [15:0] and_766__out;
  coreir_and #(.width(16)) and_766(
    .in0(and_766__in0),
    .in1(and_766__in1),
    .out(and_766__out)
  );

  //Wire declarations for instance 'and_768' (Module coreir_and)
  wire [15:0] and_768__in0;
  wire [15:0] and_768__in1;
  wire [15:0] and_768__out;
  coreir_and #(.width(16)) and_768(
    .in0(and_768__in0),
    .in1(and_768__in1),
    .out(and_768__out)
  );

  //Wire declarations for instance 'and_770' (Module coreir_and)
  wire [15:0] and_770__in0;
  wire [15:0] and_770__in1;
  wire [15:0] and_770__out;
  coreir_and #(.width(16)) and_770(
    .in0(and_770__in0),
    .in1(and_770__in1),
    .out(and_770__out)
  );

  //Wire declarations for instance 'and_772' (Module coreir_and)
  wire [15:0] and_772__in0;
  wire [15:0] and_772__in1;
  wire [15:0] and_772__out;
  coreir_and #(.width(16)) and_772(
    .in0(and_772__in0),
    .in1(and_772__in1),
    .out(and_772__out)
  );

  //Wire declarations for instance 'and_774' (Module coreir_and)
  wire [15:0] and_774__in0;
  wire [15:0] and_774__in1;
  wire [15:0] and_774__out;
  coreir_and #(.width(16)) and_774(
    .in0(and_774__in0),
    .in1(and_774__in1),
    .out(and_774__out)
  );

  //Wire declarations for instance 'and_776' (Module coreir_and)
  wire [15:0] and_776__in0;
  wire [15:0] and_776__in1;
  wire [15:0] and_776__out;
  coreir_and #(.width(16)) and_776(
    .in0(and_776__in0),
    .in1(and_776__in1),
    .out(and_776__out)
  );

  //Wire declarations for instance 'and_778' (Module coreir_and)
  wire [15:0] and_778__in0;
  wire [15:0] and_778__in1;
  wire [15:0] and_778__out;
  coreir_and #(.width(16)) and_778(
    .in0(and_778__in0),
    .in1(and_778__in1),
    .out(and_778__out)
  );

  //Wire declarations for instance 'and_78' (Module coreir_and)
  wire [15:0] and_78__in0;
  wire [15:0] and_78__in1;
  wire [15:0] and_78__out;
  coreir_and #(.width(16)) and_78(
    .in0(and_78__in0),
    .in1(and_78__in1),
    .out(and_78__out)
  );

  //Wire declarations for instance 'and_780' (Module coreir_and)
  wire [15:0] and_780__in0;
  wire [15:0] and_780__in1;
  wire [15:0] and_780__out;
  coreir_and #(.width(16)) and_780(
    .in0(and_780__in0),
    .in1(and_780__in1),
    .out(and_780__out)
  );

  //Wire declarations for instance 'and_782' (Module coreir_and)
  wire [15:0] and_782__in0;
  wire [15:0] and_782__in1;
  wire [15:0] and_782__out;
  coreir_and #(.width(16)) and_782(
    .in0(and_782__in0),
    .in1(and_782__in1),
    .out(and_782__out)
  );

  //Wire declarations for instance 'and_784' (Module coreir_and)
  wire [15:0] and_784__in0;
  wire [15:0] and_784__in1;
  wire [15:0] and_784__out;
  coreir_and #(.width(16)) and_784(
    .in0(and_784__in0),
    .in1(and_784__in1),
    .out(and_784__out)
  );

  //Wire declarations for instance 'and_786' (Module coreir_and)
  wire [15:0] and_786__in0;
  wire [15:0] and_786__in1;
  wire [15:0] and_786__out;
  coreir_and #(.width(16)) and_786(
    .in0(and_786__in0),
    .in1(and_786__in1),
    .out(and_786__out)
  );

  //Wire declarations for instance 'and_788' (Module coreir_and)
  wire [15:0] and_788__in0;
  wire [15:0] and_788__in1;
  wire [15:0] and_788__out;
  coreir_and #(.width(16)) and_788(
    .in0(and_788__in0),
    .in1(and_788__in1),
    .out(and_788__out)
  );

  //Wire declarations for instance 'and_790' (Module coreir_and)
  wire [15:0] and_790__in0;
  wire [15:0] and_790__in1;
  wire [15:0] and_790__out;
  coreir_and #(.width(16)) and_790(
    .in0(and_790__in0),
    .in1(and_790__in1),
    .out(and_790__out)
  );

  //Wire declarations for instance 'and_792' (Module coreir_and)
  wire [15:0] and_792__in0;
  wire [15:0] and_792__in1;
  wire [15:0] and_792__out;
  coreir_and #(.width(16)) and_792(
    .in0(and_792__in0),
    .in1(and_792__in1),
    .out(and_792__out)
  );

  //Wire declarations for instance 'and_794' (Module coreir_and)
  wire [15:0] and_794__in0;
  wire [15:0] and_794__in1;
  wire [15:0] and_794__out;
  coreir_and #(.width(16)) and_794(
    .in0(and_794__in0),
    .in1(and_794__in1),
    .out(and_794__out)
  );

  //Wire declarations for instance 'and_796' (Module coreir_and)
  wire [15:0] and_796__in0;
  wire [15:0] and_796__in1;
  wire [15:0] and_796__out;
  coreir_and #(.width(16)) and_796(
    .in0(and_796__in0),
    .in1(and_796__in1),
    .out(and_796__out)
  );

  //Wire declarations for instance 'and_798' (Module coreir_and)
  wire [15:0] and_798__in0;
  wire [15:0] and_798__in1;
  wire [15:0] and_798__out;
  coreir_and #(.width(16)) and_798(
    .in0(and_798__in0),
    .in1(and_798__in1),
    .out(and_798__out)
  );

  //Wire declarations for instance 'and_8' (Module coreir_and)
  wire [15:0] and_8__in0;
  wire [15:0] and_8__in1;
  wire [15:0] and_8__out;
  coreir_and #(.width(16)) and_8(
    .in0(and_8__in0),
    .in1(and_8__in1),
    .out(and_8__out)
  );

  //Wire declarations for instance 'and_80' (Module coreir_and)
  wire [15:0] and_80__in0;
  wire [15:0] and_80__in1;
  wire [15:0] and_80__out;
  coreir_and #(.width(16)) and_80(
    .in0(and_80__in0),
    .in1(and_80__in1),
    .out(and_80__out)
  );

  //Wire declarations for instance 'and_800' (Module coreir_and)
  wire [15:0] and_800__in0;
  wire [15:0] and_800__in1;
  wire [15:0] and_800__out;
  coreir_and #(.width(16)) and_800(
    .in0(and_800__in0),
    .in1(and_800__in1),
    .out(and_800__out)
  );

  //Wire declarations for instance 'and_802' (Module coreir_and)
  wire [15:0] and_802__in0;
  wire [15:0] and_802__in1;
  wire [15:0] and_802__out;
  coreir_and #(.width(16)) and_802(
    .in0(and_802__in0),
    .in1(and_802__in1),
    .out(and_802__out)
  );

  //Wire declarations for instance 'and_804' (Module coreir_and)
  wire [15:0] and_804__in0;
  wire [15:0] and_804__in1;
  wire [15:0] and_804__out;
  coreir_and #(.width(16)) and_804(
    .in0(and_804__in0),
    .in1(and_804__in1),
    .out(and_804__out)
  );

  //Wire declarations for instance 'and_806' (Module coreir_and)
  wire [15:0] and_806__in0;
  wire [15:0] and_806__in1;
  wire [15:0] and_806__out;
  coreir_and #(.width(16)) and_806(
    .in0(and_806__in0),
    .in1(and_806__in1),
    .out(and_806__out)
  );

  //Wire declarations for instance 'and_808' (Module coreir_and)
  wire [15:0] and_808__in0;
  wire [15:0] and_808__in1;
  wire [15:0] and_808__out;
  coreir_and #(.width(16)) and_808(
    .in0(and_808__in0),
    .in1(and_808__in1),
    .out(and_808__out)
  );

  //Wire declarations for instance 'and_810' (Module coreir_and)
  wire [15:0] and_810__in0;
  wire [15:0] and_810__in1;
  wire [15:0] and_810__out;
  coreir_and #(.width(16)) and_810(
    .in0(and_810__in0),
    .in1(and_810__in1),
    .out(and_810__out)
  );

  //Wire declarations for instance 'and_812' (Module coreir_and)
  wire [15:0] and_812__in0;
  wire [15:0] and_812__in1;
  wire [15:0] and_812__out;
  coreir_and #(.width(16)) and_812(
    .in0(and_812__in0),
    .in1(and_812__in1),
    .out(and_812__out)
  );

  //Wire declarations for instance 'and_814' (Module coreir_and)
  wire [15:0] and_814__in0;
  wire [15:0] and_814__in1;
  wire [15:0] and_814__out;
  coreir_and #(.width(16)) and_814(
    .in0(and_814__in0),
    .in1(and_814__in1),
    .out(and_814__out)
  );

  //Wire declarations for instance 'and_816' (Module coreir_and)
  wire [15:0] and_816__in0;
  wire [15:0] and_816__in1;
  wire [15:0] and_816__out;
  coreir_and #(.width(16)) and_816(
    .in0(and_816__in0),
    .in1(and_816__in1),
    .out(and_816__out)
  );

  //Wire declarations for instance 'and_818' (Module coreir_and)
  wire [15:0] and_818__in0;
  wire [15:0] and_818__in1;
  wire [15:0] and_818__out;
  coreir_and #(.width(16)) and_818(
    .in0(and_818__in0),
    .in1(and_818__in1),
    .out(and_818__out)
  );

  //Wire declarations for instance 'and_82' (Module coreir_and)
  wire [15:0] and_82__in0;
  wire [15:0] and_82__in1;
  wire [15:0] and_82__out;
  coreir_and #(.width(16)) and_82(
    .in0(and_82__in0),
    .in1(and_82__in1),
    .out(and_82__out)
  );

  //Wire declarations for instance 'and_820' (Module coreir_and)
  wire [15:0] and_820__in0;
  wire [15:0] and_820__in1;
  wire [15:0] and_820__out;
  coreir_and #(.width(16)) and_820(
    .in0(and_820__in0),
    .in1(and_820__in1),
    .out(and_820__out)
  );

  //Wire declarations for instance 'and_822' (Module coreir_and)
  wire [15:0] and_822__in0;
  wire [15:0] and_822__in1;
  wire [15:0] and_822__out;
  coreir_and #(.width(16)) and_822(
    .in0(and_822__in0),
    .in1(and_822__in1),
    .out(and_822__out)
  );

  //Wire declarations for instance 'and_824' (Module coreir_and)
  wire [15:0] and_824__in0;
  wire [15:0] and_824__in1;
  wire [15:0] and_824__out;
  coreir_and #(.width(16)) and_824(
    .in0(and_824__in0),
    .in1(and_824__in1),
    .out(and_824__out)
  );

  //Wire declarations for instance 'and_826' (Module coreir_and)
  wire [15:0] and_826__in0;
  wire [15:0] and_826__in1;
  wire [15:0] and_826__out;
  coreir_and #(.width(16)) and_826(
    .in0(and_826__in0),
    .in1(and_826__in1),
    .out(and_826__out)
  );

  //Wire declarations for instance 'and_828' (Module coreir_and)
  wire [15:0] and_828__in0;
  wire [15:0] and_828__in1;
  wire [15:0] and_828__out;
  coreir_and #(.width(16)) and_828(
    .in0(and_828__in0),
    .in1(and_828__in1),
    .out(and_828__out)
  );

  //Wire declarations for instance 'and_830' (Module coreir_and)
  wire [15:0] and_830__in0;
  wire [15:0] and_830__in1;
  wire [15:0] and_830__out;
  coreir_and #(.width(16)) and_830(
    .in0(and_830__in0),
    .in1(and_830__in1),
    .out(and_830__out)
  );

  //Wire declarations for instance 'and_832' (Module coreir_and)
  wire [15:0] and_832__in0;
  wire [15:0] and_832__in1;
  wire [15:0] and_832__out;
  coreir_and #(.width(16)) and_832(
    .in0(and_832__in0),
    .in1(and_832__in1),
    .out(and_832__out)
  );

  //Wire declarations for instance 'and_834' (Module coreir_and)
  wire [15:0] and_834__in0;
  wire [15:0] and_834__in1;
  wire [15:0] and_834__out;
  coreir_and #(.width(16)) and_834(
    .in0(and_834__in0),
    .in1(and_834__in1),
    .out(and_834__out)
  );

  //Wire declarations for instance 'and_836' (Module coreir_and)
  wire [15:0] and_836__in0;
  wire [15:0] and_836__in1;
  wire [15:0] and_836__out;
  coreir_and #(.width(16)) and_836(
    .in0(and_836__in0),
    .in1(and_836__in1),
    .out(and_836__out)
  );

  //Wire declarations for instance 'and_838' (Module coreir_and)
  wire [15:0] and_838__in0;
  wire [15:0] and_838__in1;
  wire [15:0] and_838__out;
  coreir_and #(.width(16)) and_838(
    .in0(and_838__in0),
    .in1(and_838__in1),
    .out(and_838__out)
  );

  //Wire declarations for instance 'and_84' (Module coreir_and)
  wire [15:0] and_84__in0;
  wire [15:0] and_84__in1;
  wire [15:0] and_84__out;
  coreir_and #(.width(16)) and_84(
    .in0(and_84__in0),
    .in1(and_84__in1),
    .out(and_84__out)
  );

  //Wire declarations for instance 'and_840' (Module coreir_and)
  wire [15:0] and_840__in0;
  wire [15:0] and_840__in1;
  wire [15:0] and_840__out;
  coreir_and #(.width(16)) and_840(
    .in0(and_840__in0),
    .in1(and_840__in1),
    .out(and_840__out)
  );

  //Wire declarations for instance 'and_842' (Module coreir_and)
  wire [15:0] and_842__in0;
  wire [15:0] and_842__in1;
  wire [15:0] and_842__out;
  coreir_and #(.width(16)) and_842(
    .in0(and_842__in0),
    .in1(and_842__in1),
    .out(and_842__out)
  );

  //Wire declarations for instance 'and_844' (Module coreir_and)
  wire [15:0] and_844__in0;
  wire [15:0] and_844__in1;
  wire [15:0] and_844__out;
  coreir_and #(.width(16)) and_844(
    .in0(and_844__in0),
    .in1(and_844__in1),
    .out(and_844__out)
  );

  //Wire declarations for instance 'and_846' (Module coreir_and)
  wire [15:0] and_846__in0;
  wire [15:0] and_846__in1;
  wire [15:0] and_846__out;
  coreir_and #(.width(16)) and_846(
    .in0(and_846__in0),
    .in1(and_846__in1),
    .out(and_846__out)
  );

  //Wire declarations for instance 'and_848' (Module coreir_and)
  wire [15:0] and_848__in0;
  wire [15:0] and_848__in1;
  wire [15:0] and_848__out;
  coreir_and #(.width(16)) and_848(
    .in0(and_848__in0),
    .in1(and_848__in1),
    .out(and_848__out)
  );

  //Wire declarations for instance 'and_850' (Module coreir_and)
  wire [15:0] and_850__in0;
  wire [15:0] and_850__in1;
  wire [15:0] and_850__out;
  coreir_and #(.width(16)) and_850(
    .in0(and_850__in0),
    .in1(and_850__in1),
    .out(and_850__out)
  );

  //Wire declarations for instance 'and_852' (Module coreir_and)
  wire [15:0] and_852__in0;
  wire [15:0] and_852__in1;
  wire [15:0] and_852__out;
  coreir_and #(.width(16)) and_852(
    .in0(and_852__in0),
    .in1(and_852__in1),
    .out(and_852__out)
  );

  //Wire declarations for instance 'and_854' (Module coreir_and)
  wire [15:0] and_854__in0;
  wire [15:0] and_854__in1;
  wire [15:0] and_854__out;
  coreir_and #(.width(16)) and_854(
    .in0(and_854__in0),
    .in1(and_854__in1),
    .out(and_854__out)
  );

  //Wire declarations for instance 'and_856' (Module coreir_and)
  wire [15:0] and_856__in0;
  wire [15:0] and_856__in1;
  wire [15:0] and_856__out;
  coreir_and #(.width(16)) and_856(
    .in0(and_856__in0),
    .in1(and_856__in1),
    .out(and_856__out)
  );

  //Wire declarations for instance 'and_858' (Module coreir_and)
  wire [15:0] and_858__in0;
  wire [15:0] and_858__in1;
  wire [15:0] and_858__out;
  coreir_and #(.width(16)) and_858(
    .in0(and_858__in0),
    .in1(and_858__in1),
    .out(and_858__out)
  );

  //Wire declarations for instance 'and_86' (Module coreir_and)
  wire [15:0] and_86__in0;
  wire [15:0] and_86__in1;
  wire [15:0] and_86__out;
  coreir_and #(.width(16)) and_86(
    .in0(and_86__in0),
    .in1(and_86__in1),
    .out(and_86__out)
  );

  //Wire declarations for instance 'and_860' (Module coreir_and)
  wire [15:0] and_860__in0;
  wire [15:0] and_860__in1;
  wire [15:0] and_860__out;
  coreir_and #(.width(16)) and_860(
    .in0(and_860__in0),
    .in1(and_860__in1),
    .out(and_860__out)
  );

  //Wire declarations for instance 'and_862' (Module coreir_and)
  wire [15:0] and_862__in0;
  wire [15:0] and_862__in1;
  wire [15:0] and_862__out;
  coreir_and #(.width(16)) and_862(
    .in0(and_862__in0),
    .in1(and_862__in1),
    .out(and_862__out)
  );

  //Wire declarations for instance 'and_864' (Module coreir_and)
  wire [15:0] and_864__in0;
  wire [15:0] and_864__in1;
  wire [15:0] and_864__out;
  coreir_and #(.width(16)) and_864(
    .in0(and_864__in0),
    .in1(and_864__in1),
    .out(and_864__out)
  );

  //Wire declarations for instance 'and_866' (Module coreir_and)
  wire [15:0] and_866__in0;
  wire [15:0] and_866__in1;
  wire [15:0] and_866__out;
  coreir_and #(.width(16)) and_866(
    .in0(and_866__in0),
    .in1(and_866__in1),
    .out(and_866__out)
  );

  //Wire declarations for instance 'and_868' (Module coreir_and)
  wire [15:0] and_868__in0;
  wire [15:0] and_868__in1;
  wire [15:0] and_868__out;
  coreir_and #(.width(16)) and_868(
    .in0(and_868__in0),
    .in1(and_868__in1),
    .out(and_868__out)
  );

  //Wire declarations for instance 'and_870' (Module coreir_and)
  wire [15:0] and_870__in0;
  wire [15:0] and_870__in1;
  wire [15:0] and_870__out;
  coreir_and #(.width(16)) and_870(
    .in0(and_870__in0),
    .in1(and_870__in1),
    .out(and_870__out)
  );

  //Wire declarations for instance 'and_872' (Module coreir_and)
  wire [15:0] and_872__in0;
  wire [15:0] and_872__in1;
  wire [15:0] and_872__out;
  coreir_and #(.width(16)) and_872(
    .in0(and_872__in0),
    .in1(and_872__in1),
    .out(and_872__out)
  );

  //Wire declarations for instance 'and_874' (Module coreir_and)
  wire [15:0] and_874__in0;
  wire [15:0] and_874__in1;
  wire [15:0] and_874__out;
  coreir_and #(.width(16)) and_874(
    .in0(and_874__in0),
    .in1(and_874__in1),
    .out(and_874__out)
  );

  //Wire declarations for instance 'and_876' (Module coreir_and)
  wire [15:0] and_876__in0;
  wire [15:0] and_876__in1;
  wire [15:0] and_876__out;
  coreir_and #(.width(16)) and_876(
    .in0(and_876__in0),
    .in1(and_876__in1),
    .out(and_876__out)
  );

  //Wire declarations for instance 'and_878' (Module coreir_and)
  wire [15:0] and_878__in0;
  wire [15:0] and_878__in1;
  wire [15:0] and_878__out;
  coreir_and #(.width(16)) and_878(
    .in0(and_878__in0),
    .in1(and_878__in1),
    .out(and_878__out)
  );

  //Wire declarations for instance 'and_88' (Module coreir_and)
  wire [15:0] and_88__in0;
  wire [15:0] and_88__in1;
  wire [15:0] and_88__out;
  coreir_and #(.width(16)) and_88(
    .in0(and_88__in0),
    .in1(and_88__in1),
    .out(and_88__out)
  );

  //Wire declarations for instance 'and_880' (Module coreir_and)
  wire [15:0] and_880__in0;
  wire [15:0] and_880__in1;
  wire [15:0] and_880__out;
  coreir_and #(.width(16)) and_880(
    .in0(and_880__in0),
    .in1(and_880__in1),
    .out(and_880__out)
  );

  //Wire declarations for instance 'and_882' (Module coreir_and)
  wire [15:0] and_882__in0;
  wire [15:0] and_882__in1;
  wire [15:0] and_882__out;
  coreir_and #(.width(16)) and_882(
    .in0(and_882__in0),
    .in1(and_882__in1),
    .out(and_882__out)
  );

  //Wire declarations for instance 'and_884' (Module coreir_and)
  wire [15:0] and_884__in0;
  wire [15:0] and_884__in1;
  wire [15:0] and_884__out;
  coreir_and #(.width(16)) and_884(
    .in0(and_884__in0),
    .in1(and_884__in1),
    .out(and_884__out)
  );

  //Wire declarations for instance 'and_886' (Module coreir_and)
  wire [15:0] and_886__in0;
  wire [15:0] and_886__in1;
  wire [15:0] and_886__out;
  coreir_and #(.width(16)) and_886(
    .in0(and_886__in0),
    .in1(and_886__in1),
    .out(and_886__out)
  );

  //Wire declarations for instance 'and_888' (Module coreir_and)
  wire [15:0] and_888__in0;
  wire [15:0] and_888__in1;
  wire [15:0] and_888__out;
  coreir_and #(.width(16)) and_888(
    .in0(and_888__in0),
    .in1(and_888__in1),
    .out(and_888__out)
  );

  //Wire declarations for instance 'and_890' (Module coreir_and)
  wire [15:0] and_890__in0;
  wire [15:0] and_890__in1;
  wire [15:0] and_890__out;
  coreir_and #(.width(16)) and_890(
    .in0(and_890__in0),
    .in1(and_890__in1),
    .out(and_890__out)
  );

  //Wire declarations for instance 'and_892' (Module coreir_and)
  wire [15:0] and_892__in0;
  wire [15:0] and_892__in1;
  wire [15:0] and_892__out;
  coreir_and #(.width(16)) and_892(
    .in0(and_892__in0),
    .in1(and_892__in1),
    .out(and_892__out)
  );

  //Wire declarations for instance 'and_894' (Module coreir_and)
  wire [15:0] and_894__in0;
  wire [15:0] and_894__in1;
  wire [15:0] and_894__out;
  coreir_and #(.width(16)) and_894(
    .in0(and_894__in0),
    .in1(and_894__in1),
    .out(and_894__out)
  );

  //Wire declarations for instance 'and_896' (Module coreir_and)
  wire [15:0] and_896__in0;
  wire [15:0] and_896__in1;
  wire [15:0] and_896__out;
  coreir_and #(.width(16)) and_896(
    .in0(and_896__in0),
    .in1(and_896__in1),
    .out(and_896__out)
  );

  //Wire declarations for instance 'and_898' (Module coreir_and)
  wire [15:0] and_898__in0;
  wire [15:0] and_898__in1;
  wire [15:0] and_898__out;
  coreir_and #(.width(16)) and_898(
    .in0(and_898__in0),
    .in1(and_898__in1),
    .out(and_898__out)
  );

  //Wire declarations for instance 'and_90' (Module coreir_and)
  wire [15:0] and_90__in0;
  wire [15:0] and_90__in1;
  wire [15:0] and_90__out;
  coreir_and #(.width(16)) and_90(
    .in0(and_90__in0),
    .in1(and_90__in1),
    .out(and_90__out)
  );

  //Wire declarations for instance 'and_900' (Module coreir_and)
  wire [15:0] and_900__in0;
  wire [15:0] and_900__in1;
  wire [15:0] and_900__out;
  coreir_and #(.width(16)) and_900(
    .in0(and_900__in0),
    .in1(and_900__in1),
    .out(and_900__out)
  );

  //Wire declarations for instance 'and_902' (Module coreir_and)
  wire [15:0] and_902__in0;
  wire [15:0] and_902__in1;
  wire [15:0] and_902__out;
  coreir_and #(.width(16)) and_902(
    .in0(and_902__in0),
    .in1(and_902__in1),
    .out(and_902__out)
  );

  //Wire declarations for instance 'and_904' (Module coreir_and)
  wire [15:0] and_904__in0;
  wire [15:0] and_904__in1;
  wire [15:0] and_904__out;
  coreir_and #(.width(16)) and_904(
    .in0(and_904__in0),
    .in1(and_904__in1),
    .out(and_904__out)
  );

  //Wire declarations for instance 'and_906' (Module coreir_and)
  wire [15:0] and_906__in0;
  wire [15:0] and_906__in1;
  wire [15:0] and_906__out;
  coreir_and #(.width(16)) and_906(
    .in0(and_906__in0),
    .in1(and_906__in1),
    .out(and_906__out)
  );

  //Wire declarations for instance 'and_908' (Module coreir_and)
  wire [15:0] and_908__in0;
  wire [15:0] and_908__in1;
  wire [15:0] and_908__out;
  coreir_and #(.width(16)) and_908(
    .in0(and_908__in0),
    .in1(and_908__in1),
    .out(and_908__out)
  );

  //Wire declarations for instance 'and_910' (Module coreir_and)
  wire [15:0] and_910__in0;
  wire [15:0] and_910__in1;
  wire [15:0] and_910__out;
  coreir_and #(.width(16)) and_910(
    .in0(and_910__in0),
    .in1(and_910__in1),
    .out(and_910__out)
  );

  //Wire declarations for instance 'and_912' (Module coreir_and)
  wire [15:0] and_912__in0;
  wire [15:0] and_912__in1;
  wire [15:0] and_912__out;
  coreir_and #(.width(16)) and_912(
    .in0(and_912__in0),
    .in1(and_912__in1),
    .out(and_912__out)
  );

  //Wire declarations for instance 'and_914' (Module coreir_and)
  wire [15:0] and_914__in0;
  wire [15:0] and_914__in1;
  wire [15:0] and_914__out;
  coreir_and #(.width(16)) and_914(
    .in0(and_914__in0),
    .in1(and_914__in1),
    .out(and_914__out)
  );

  //Wire declarations for instance 'and_916' (Module coreir_and)
  wire [15:0] and_916__in0;
  wire [15:0] and_916__in1;
  wire [15:0] and_916__out;
  coreir_and #(.width(16)) and_916(
    .in0(and_916__in0),
    .in1(and_916__in1),
    .out(and_916__out)
  );

  //Wire declarations for instance 'and_918' (Module coreir_and)
  wire [15:0] and_918__in0;
  wire [15:0] and_918__in1;
  wire [15:0] and_918__out;
  coreir_and #(.width(16)) and_918(
    .in0(and_918__in0),
    .in1(and_918__in1),
    .out(and_918__out)
  );

  //Wire declarations for instance 'and_92' (Module coreir_and)
  wire [15:0] and_92__in0;
  wire [15:0] and_92__in1;
  wire [15:0] and_92__out;
  coreir_and #(.width(16)) and_92(
    .in0(and_92__in0),
    .in1(and_92__in1),
    .out(and_92__out)
  );

  //Wire declarations for instance 'and_920' (Module coreir_and)
  wire [15:0] and_920__in0;
  wire [15:0] and_920__in1;
  wire [15:0] and_920__out;
  coreir_and #(.width(16)) and_920(
    .in0(and_920__in0),
    .in1(and_920__in1),
    .out(and_920__out)
  );

  //Wire declarations for instance 'and_922' (Module coreir_and)
  wire [15:0] and_922__in0;
  wire [15:0] and_922__in1;
  wire [15:0] and_922__out;
  coreir_and #(.width(16)) and_922(
    .in0(and_922__in0),
    .in1(and_922__in1),
    .out(and_922__out)
  );

  //Wire declarations for instance 'and_924' (Module coreir_and)
  wire [15:0] and_924__in0;
  wire [15:0] and_924__in1;
  wire [15:0] and_924__out;
  coreir_and #(.width(16)) and_924(
    .in0(and_924__in0),
    .in1(and_924__in1),
    .out(and_924__out)
  );

  //Wire declarations for instance 'and_926' (Module coreir_and)
  wire [15:0] and_926__in0;
  wire [15:0] and_926__in1;
  wire [15:0] and_926__out;
  coreir_and #(.width(16)) and_926(
    .in0(and_926__in0),
    .in1(and_926__in1),
    .out(and_926__out)
  );

  //Wire declarations for instance 'and_928' (Module coreir_and)
  wire [15:0] and_928__in0;
  wire [15:0] and_928__in1;
  wire [15:0] and_928__out;
  coreir_and #(.width(16)) and_928(
    .in0(and_928__in0),
    .in1(and_928__in1),
    .out(and_928__out)
  );

  //Wire declarations for instance 'and_930' (Module coreir_and)
  wire [15:0] and_930__in0;
  wire [15:0] and_930__in1;
  wire [15:0] and_930__out;
  coreir_and #(.width(16)) and_930(
    .in0(and_930__in0),
    .in1(and_930__in1),
    .out(and_930__out)
  );

  //Wire declarations for instance 'and_932' (Module coreir_and)
  wire [15:0] and_932__in0;
  wire [15:0] and_932__in1;
  wire [15:0] and_932__out;
  coreir_and #(.width(16)) and_932(
    .in0(and_932__in0),
    .in1(and_932__in1),
    .out(and_932__out)
  );

  //Wire declarations for instance 'and_934' (Module coreir_and)
  wire [15:0] and_934__in0;
  wire [15:0] and_934__in1;
  wire [15:0] and_934__out;
  coreir_and #(.width(16)) and_934(
    .in0(and_934__in0),
    .in1(and_934__in1),
    .out(and_934__out)
  );

  //Wire declarations for instance 'and_936' (Module coreir_and)
  wire [15:0] and_936__in0;
  wire [15:0] and_936__in1;
  wire [15:0] and_936__out;
  coreir_and #(.width(16)) and_936(
    .in0(and_936__in0),
    .in1(and_936__in1),
    .out(and_936__out)
  );

  //Wire declarations for instance 'and_938' (Module coreir_and)
  wire [15:0] and_938__in0;
  wire [15:0] and_938__in1;
  wire [15:0] and_938__out;
  coreir_and #(.width(16)) and_938(
    .in0(and_938__in0),
    .in1(and_938__in1),
    .out(and_938__out)
  );

  //Wire declarations for instance 'and_94' (Module coreir_and)
  wire [15:0] and_94__in0;
  wire [15:0] and_94__in1;
  wire [15:0] and_94__out;
  coreir_and #(.width(16)) and_94(
    .in0(and_94__in0),
    .in1(and_94__in1),
    .out(and_94__out)
  );

  //Wire declarations for instance 'and_940' (Module coreir_and)
  wire [15:0] and_940__in0;
  wire [15:0] and_940__in1;
  wire [15:0] and_940__out;
  coreir_and #(.width(16)) and_940(
    .in0(and_940__in0),
    .in1(and_940__in1),
    .out(and_940__out)
  );

  //Wire declarations for instance 'and_942' (Module coreir_and)
  wire [15:0] and_942__in0;
  wire [15:0] and_942__in1;
  wire [15:0] and_942__out;
  coreir_and #(.width(16)) and_942(
    .in0(and_942__in0),
    .in1(and_942__in1),
    .out(and_942__out)
  );

  //Wire declarations for instance 'and_944' (Module coreir_and)
  wire [15:0] and_944__in0;
  wire [15:0] and_944__in1;
  wire [15:0] and_944__out;
  coreir_and #(.width(16)) and_944(
    .in0(and_944__in0),
    .in1(and_944__in1),
    .out(and_944__out)
  );

  //Wire declarations for instance 'and_946' (Module coreir_and)
  wire [15:0] and_946__in0;
  wire [15:0] and_946__in1;
  wire [15:0] and_946__out;
  coreir_and #(.width(16)) and_946(
    .in0(and_946__in0),
    .in1(and_946__in1),
    .out(and_946__out)
  );

  //Wire declarations for instance 'and_948' (Module coreir_and)
  wire [15:0] and_948__in0;
  wire [15:0] and_948__in1;
  wire [15:0] and_948__out;
  coreir_and #(.width(16)) and_948(
    .in0(and_948__in0),
    .in1(and_948__in1),
    .out(and_948__out)
  );

  //Wire declarations for instance 'and_950' (Module coreir_and)
  wire [15:0] and_950__in0;
  wire [15:0] and_950__in1;
  wire [15:0] and_950__out;
  coreir_and #(.width(16)) and_950(
    .in0(and_950__in0),
    .in1(and_950__in1),
    .out(and_950__out)
  );

  //Wire declarations for instance 'and_952' (Module coreir_and)
  wire [15:0] and_952__in0;
  wire [15:0] and_952__in1;
  wire [15:0] and_952__out;
  coreir_and #(.width(16)) and_952(
    .in0(and_952__in0),
    .in1(and_952__in1),
    .out(and_952__out)
  );

  //Wire declarations for instance 'and_954' (Module coreir_and)
  wire [15:0] and_954__in0;
  wire [15:0] and_954__in1;
  wire [15:0] and_954__out;
  coreir_and #(.width(16)) and_954(
    .in0(and_954__in0),
    .in1(and_954__in1),
    .out(and_954__out)
  );

  //Wire declarations for instance 'and_956' (Module coreir_and)
  wire [15:0] and_956__in0;
  wire [15:0] and_956__in1;
  wire [15:0] and_956__out;
  coreir_and #(.width(16)) and_956(
    .in0(and_956__in0),
    .in1(and_956__in1),
    .out(and_956__out)
  );

  //Wire declarations for instance 'and_958' (Module coreir_and)
  wire [15:0] and_958__in0;
  wire [15:0] and_958__in1;
  wire [15:0] and_958__out;
  coreir_and #(.width(16)) and_958(
    .in0(and_958__in0),
    .in1(and_958__in1),
    .out(and_958__out)
  );

  //Wire declarations for instance 'and_96' (Module coreir_and)
  wire [15:0] and_96__in0;
  wire [15:0] and_96__in1;
  wire [15:0] and_96__out;
  coreir_and #(.width(16)) and_96(
    .in0(and_96__in0),
    .in1(and_96__in1),
    .out(and_96__out)
  );

  //Wire declarations for instance 'and_960' (Module coreir_and)
  wire [15:0] and_960__in0;
  wire [15:0] and_960__in1;
  wire [15:0] and_960__out;
  coreir_and #(.width(16)) and_960(
    .in0(and_960__in0),
    .in1(and_960__in1),
    .out(and_960__out)
  );

  //Wire declarations for instance 'and_962' (Module coreir_and)
  wire [15:0] and_962__in0;
  wire [15:0] and_962__in1;
  wire [15:0] and_962__out;
  coreir_and #(.width(16)) and_962(
    .in0(and_962__in0),
    .in1(and_962__in1),
    .out(and_962__out)
  );

  //Wire declarations for instance 'and_964' (Module coreir_and)
  wire [15:0] and_964__in0;
  wire [15:0] and_964__in1;
  wire [15:0] and_964__out;
  coreir_and #(.width(16)) and_964(
    .in0(and_964__in0),
    .in1(and_964__in1),
    .out(and_964__out)
  );

  //Wire declarations for instance 'and_966' (Module coreir_and)
  wire [15:0] and_966__in0;
  wire [15:0] and_966__in1;
  wire [15:0] and_966__out;
  coreir_and #(.width(16)) and_966(
    .in0(and_966__in0),
    .in1(and_966__in1),
    .out(and_966__out)
  );

  //Wire declarations for instance 'and_968' (Module coreir_and)
  wire [15:0] and_968__in0;
  wire [15:0] and_968__in1;
  wire [15:0] and_968__out;
  coreir_and #(.width(16)) and_968(
    .in0(and_968__in0),
    .in1(and_968__in1),
    .out(and_968__out)
  );

  //Wire declarations for instance 'and_970' (Module coreir_and)
  wire [15:0] and_970__in0;
  wire [15:0] and_970__in1;
  wire [15:0] and_970__out;
  coreir_and #(.width(16)) and_970(
    .in0(and_970__in0),
    .in1(and_970__in1),
    .out(and_970__out)
  );

  //Wire declarations for instance 'and_972' (Module coreir_and)
  wire [15:0] and_972__in0;
  wire [15:0] and_972__in1;
  wire [15:0] and_972__out;
  coreir_and #(.width(16)) and_972(
    .in0(and_972__in0),
    .in1(and_972__in1),
    .out(and_972__out)
  );

  //Wire declarations for instance 'and_974' (Module coreir_and)
  wire [15:0] and_974__in0;
  wire [15:0] and_974__in1;
  wire [15:0] and_974__out;
  coreir_and #(.width(16)) and_974(
    .in0(and_974__in0),
    .in1(and_974__in1),
    .out(and_974__out)
  );

  //Wire declarations for instance 'and_976' (Module coreir_and)
  wire [15:0] and_976__in0;
  wire [15:0] and_976__in1;
  wire [15:0] and_976__out;
  coreir_and #(.width(16)) and_976(
    .in0(and_976__in0),
    .in1(and_976__in1),
    .out(and_976__out)
  );

  //Wire declarations for instance 'and_978' (Module coreir_and)
  wire [15:0] and_978__in0;
  wire [15:0] and_978__in1;
  wire [15:0] and_978__out;
  coreir_and #(.width(16)) and_978(
    .in0(and_978__in0),
    .in1(and_978__in1),
    .out(and_978__out)
  );

  //Wire declarations for instance 'and_98' (Module coreir_and)
  wire [15:0] and_98__in0;
  wire [15:0] and_98__in1;
  wire [15:0] and_98__out;
  coreir_and #(.width(16)) and_98(
    .in0(and_98__in0),
    .in1(and_98__in1),
    .out(and_98__out)
  );

  //Wire declarations for instance 'and_980' (Module coreir_and)
  wire [15:0] and_980__in0;
  wire [15:0] and_980__in1;
  wire [15:0] and_980__out;
  coreir_and #(.width(16)) and_980(
    .in0(and_980__in0),
    .in1(and_980__in1),
    .out(and_980__out)
  );

  //Wire declarations for instance 'and_982' (Module coreir_and)
  wire [15:0] and_982__in0;
  wire [15:0] and_982__in1;
  wire [15:0] and_982__out;
  coreir_and #(.width(16)) and_982(
    .in0(and_982__in0),
    .in1(and_982__in1),
    .out(and_982__out)
  );

  //Wire declarations for instance 'and_984' (Module coreir_and)
  wire [15:0] and_984__in0;
  wire [15:0] and_984__in1;
  wire [15:0] and_984__out;
  coreir_and #(.width(16)) and_984(
    .in0(and_984__in0),
    .in1(and_984__in1),
    .out(and_984__out)
  );

  //Wire declarations for instance 'and_986' (Module coreir_and)
  wire [15:0] and_986__in0;
  wire [15:0] and_986__in1;
  wire [15:0] and_986__out;
  coreir_and #(.width(16)) and_986(
    .in0(and_986__in0),
    .in1(and_986__in1),
    .out(and_986__out)
  );

  //Wire declarations for instance 'and_988' (Module coreir_and)
  wire [15:0] and_988__in0;
  wire [15:0] and_988__in1;
  wire [15:0] and_988__out;
  coreir_and #(.width(16)) and_988(
    .in0(and_988__in0),
    .in1(and_988__in1),
    .out(and_988__out)
  );

  //Wire declarations for instance 'and_990' (Module coreir_and)
  wire [15:0] and_990__in0;
  wire [15:0] and_990__in1;
  wire [15:0] and_990__out;
  coreir_and #(.width(16)) and_990(
    .in0(and_990__in0),
    .in1(and_990__in1),
    .out(and_990__out)
  );

  //Wire declarations for instance 'and_992' (Module coreir_and)
  wire [15:0] and_992__in0;
  wire [15:0] and_992__in1;
  wire [15:0] and_992__out;
  coreir_and #(.width(16)) and_992(
    .in0(and_992__in0),
    .in1(and_992__in1),
    .out(and_992__out)
  );

  //Wire declarations for instance 'and_994' (Module coreir_and)
  wire [15:0] and_994__in0;
  wire [15:0] and_994__in1;
  wire [15:0] and_994__out;
  coreir_and #(.width(16)) and_994(
    .in0(and_994__in0),
    .in1(and_994__in1),
    .out(and_994__out)
  );

  //Wire declarations for instance 'and_996' (Module coreir_and)
  wire [15:0] and_996__in0;
  wire [15:0] and_996__in1;
  wire [15:0] and_996__out;
  coreir_and #(.width(16)) and_996(
    .in0(and_996__in0),
    .in1(and_996__in1),
    .out(and_996__out)
  );

  //Wire declarations for instance 'and_998' (Module coreir_and)
  wire [15:0] and_998__in0;
  wire [15:0] and_998__in1;
  wire [15:0] and_998__out;
  coreir_and #(.width(16)) and_998(
    .in0(and_998__in0),
    .in1(and_998__in1),
    .out(and_998__out)
  );

  //Wire declarations for instance 'or_1' (Module coreir_or)
  wire [15:0] or_1__in0;
  wire [15:0] or_1__in1;
  wire [15:0] or_1__out;
  coreir_or #(.width(16)) or_1(
    .in0(or_1__in0),
    .in1(or_1__in1),
    .out(or_1__out)
  );

  //Wire declarations for instance 'or_101' (Module coreir_or)
  wire [15:0] or_101__in0;
  wire [15:0] or_101__in1;
  wire [15:0] or_101__out;
  coreir_or #(.width(16)) or_101(
    .in0(or_101__in0),
    .in1(or_101__in1),
    .out(or_101__out)
  );

  //Wire declarations for instance 'or_103' (Module coreir_or)
  wire [15:0] or_103__in0;
  wire [15:0] or_103__in1;
  wire [15:0] or_103__out;
  coreir_or #(.width(16)) or_103(
    .in0(or_103__in0),
    .in1(or_103__in1),
    .out(or_103__out)
  );

  //Wire declarations for instance 'or_105' (Module coreir_or)
  wire [15:0] or_105__in0;
  wire [15:0] or_105__in1;
  wire [15:0] or_105__out;
  coreir_or #(.width(16)) or_105(
    .in0(or_105__in0),
    .in1(or_105__in1),
    .out(or_105__out)
  );

  //Wire declarations for instance 'or_107' (Module coreir_or)
  wire [15:0] or_107__in0;
  wire [15:0] or_107__in1;
  wire [15:0] or_107__out;
  coreir_or #(.width(16)) or_107(
    .in0(or_107__in0),
    .in1(or_107__in1),
    .out(or_107__out)
  );

  //Wire declarations for instance 'or_109' (Module coreir_or)
  wire [15:0] or_109__in0;
  wire [15:0] or_109__in1;
  wire [15:0] or_109__out;
  coreir_or #(.width(16)) or_109(
    .in0(or_109__in0),
    .in1(or_109__in1),
    .out(or_109__out)
  );

  //Wire declarations for instance 'or_11' (Module coreir_or)
  wire [15:0] or_11__in0;
  wire [15:0] or_11__in1;
  wire [15:0] or_11__out;
  coreir_or #(.width(16)) or_11(
    .in0(or_11__in0),
    .in1(or_11__in1),
    .out(or_11__out)
  );

  //Wire declarations for instance 'or_111' (Module coreir_or)
  wire [15:0] or_111__in0;
  wire [15:0] or_111__in1;
  wire [15:0] or_111__out;
  coreir_or #(.width(16)) or_111(
    .in0(or_111__in0),
    .in1(or_111__in1),
    .out(or_111__out)
  );

  //Wire declarations for instance 'or_113' (Module coreir_or)
  wire [15:0] or_113__in0;
  wire [15:0] or_113__in1;
  wire [15:0] or_113__out;
  coreir_or #(.width(16)) or_113(
    .in0(or_113__in0),
    .in1(or_113__in1),
    .out(or_113__out)
  );

  //Wire declarations for instance 'or_115' (Module coreir_or)
  wire [15:0] or_115__in0;
  wire [15:0] or_115__in1;
  wire [15:0] or_115__out;
  coreir_or #(.width(16)) or_115(
    .in0(or_115__in0),
    .in1(or_115__in1),
    .out(or_115__out)
  );

  //Wire declarations for instance 'or_117' (Module coreir_or)
  wire [15:0] or_117__in0;
  wire [15:0] or_117__in1;
  wire [15:0] or_117__out;
  coreir_or #(.width(16)) or_117(
    .in0(or_117__in0),
    .in1(or_117__in1),
    .out(or_117__out)
  );

  //Wire declarations for instance 'or_119' (Module coreir_or)
  wire [15:0] or_119__in0;
  wire [15:0] or_119__in1;
  wire [15:0] or_119__out;
  coreir_or #(.width(16)) or_119(
    .in0(or_119__in0),
    .in1(or_119__in1),
    .out(or_119__out)
  );

  //Wire declarations for instance 'or_121' (Module coreir_or)
  wire [15:0] or_121__in0;
  wire [15:0] or_121__in1;
  wire [15:0] or_121__out;
  coreir_or #(.width(16)) or_121(
    .in0(or_121__in0),
    .in1(or_121__in1),
    .out(or_121__out)
  );

  //Wire declarations for instance 'or_123' (Module coreir_or)
  wire [15:0] or_123__in0;
  wire [15:0] or_123__in1;
  wire [15:0] or_123__out;
  coreir_or #(.width(16)) or_123(
    .in0(or_123__in0),
    .in1(or_123__in1),
    .out(or_123__out)
  );

  //Wire declarations for instance 'or_125' (Module coreir_or)
  wire [15:0] or_125__in0;
  wire [15:0] or_125__in1;
  wire [15:0] or_125__out;
  coreir_or #(.width(16)) or_125(
    .in0(or_125__in0),
    .in1(or_125__in1),
    .out(or_125__out)
  );

  //Wire declarations for instance 'or_127' (Module coreir_or)
  wire [15:0] or_127__in0;
  wire [15:0] or_127__in1;
  wire [15:0] or_127__out;
  coreir_or #(.width(16)) or_127(
    .in0(or_127__in0),
    .in1(or_127__in1),
    .out(or_127__out)
  );

  //Wire declarations for instance 'or_129' (Module coreir_or)
  wire [15:0] or_129__in0;
  wire [15:0] or_129__in1;
  wire [15:0] or_129__out;
  coreir_or #(.width(16)) or_129(
    .in0(or_129__in0),
    .in1(or_129__in1),
    .out(or_129__out)
  );

  //Wire declarations for instance 'or_13' (Module coreir_or)
  wire [15:0] or_13__in0;
  wire [15:0] or_13__in1;
  wire [15:0] or_13__out;
  coreir_or #(.width(16)) or_13(
    .in0(or_13__in0),
    .in1(or_13__in1),
    .out(or_13__out)
  );

  //Wire declarations for instance 'or_131' (Module coreir_or)
  wire [15:0] or_131__in0;
  wire [15:0] or_131__in1;
  wire [15:0] or_131__out;
  coreir_or #(.width(16)) or_131(
    .in0(or_131__in0),
    .in1(or_131__in1),
    .out(or_131__out)
  );

  //Wire declarations for instance 'or_133' (Module coreir_or)
  wire [15:0] or_133__in0;
  wire [15:0] or_133__in1;
  wire [15:0] or_133__out;
  coreir_or #(.width(16)) or_133(
    .in0(or_133__in0),
    .in1(or_133__in1),
    .out(or_133__out)
  );

  //Wire declarations for instance 'or_135' (Module coreir_or)
  wire [15:0] or_135__in0;
  wire [15:0] or_135__in1;
  wire [15:0] or_135__out;
  coreir_or #(.width(16)) or_135(
    .in0(or_135__in0),
    .in1(or_135__in1),
    .out(or_135__out)
  );

  //Wire declarations for instance 'or_137' (Module coreir_or)
  wire [15:0] or_137__in0;
  wire [15:0] or_137__in1;
  wire [15:0] or_137__out;
  coreir_or #(.width(16)) or_137(
    .in0(or_137__in0),
    .in1(or_137__in1),
    .out(or_137__out)
  );

  //Wire declarations for instance 'or_139' (Module coreir_or)
  wire [15:0] or_139__in0;
  wire [15:0] or_139__in1;
  wire [15:0] or_139__out;
  coreir_or #(.width(16)) or_139(
    .in0(or_139__in0),
    .in1(or_139__in1),
    .out(or_139__out)
  );

  //Wire declarations for instance 'or_141' (Module coreir_or)
  wire [15:0] or_141__in0;
  wire [15:0] or_141__in1;
  wire [15:0] or_141__out;
  coreir_or #(.width(16)) or_141(
    .in0(or_141__in0),
    .in1(or_141__in1),
    .out(or_141__out)
  );

  //Wire declarations for instance 'or_143' (Module coreir_or)
  wire [15:0] or_143__in0;
  wire [15:0] or_143__in1;
  wire [15:0] or_143__out;
  coreir_or #(.width(16)) or_143(
    .in0(or_143__in0),
    .in1(or_143__in1),
    .out(or_143__out)
  );

  //Wire declarations for instance 'or_145' (Module coreir_or)
  wire [15:0] or_145__in0;
  wire [15:0] or_145__in1;
  wire [15:0] or_145__out;
  coreir_or #(.width(16)) or_145(
    .in0(or_145__in0),
    .in1(or_145__in1),
    .out(or_145__out)
  );

  //Wire declarations for instance 'or_147' (Module coreir_or)
  wire [15:0] or_147__in0;
  wire [15:0] or_147__in1;
  wire [15:0] or_147__out;
  coreir_or #(.width(16)) or_147(
    .in0(or_147__in0),
    .in1(or_147__in1),
    .out(or_147__out)
  );

  //Wire declarations for instance 'or_149' (Module coreir_or)
  wire [15:0] or_149__in0;
  wire [15:0] or_149__in1;
  wire [15:0] or_149__out;
  coreir_or #(.width(16)) or_149(
    .in0(or_149__in0),
    .in1(or_149__in1),
    .out(or_149__out)
  );

  //Wire declarations for instance 'or_15' (Module coreir_or)
  wire [15:0] or_15__in0;
  wire [15:0] or_15__in1;
  wire [15:0] or_15__out;
  coreir_or #(.width(16)) or_15(
    .in0(or_15__in0),
    .in1(or_15__in1),
    .out(or_15__out)
  );

  //Wire declarations for instance 'or_151' (Module coreir_or)
  wire [15:0] or_151__in0;
  wire [15:0] or_151__in1;
  wire [15:0] or_151__out;
  coreir_or #(.width(16)) or_151(
    .in0(or_151__in0),
    .in1(or_151__in1),
    .out(or_151__out)
  );

  //Wire declarations for instance 'or_153' (Module coreir_or)
  wire [15:0] or_153__in0;
  wire [15:0] or_153__in1;
  wire [15:0] or_153__out;
  coreir_or #(.width(16)) or_153(
    .in0(or_153__in0),
    .in1(or_153__in1),
    .out(or_153__out)
  );

  //Wire declarations for instance 'or_155' (Module coreir_or)
  wire [15:0] or_155__in0;
  wire [15:0] or_155__in1;
  wire [15:0] or_155__out;
  coreir_or #(.width(16)) or_155(
    .in0(or_155__in0),
    .in1(or_155__in1),
    .out(or_155__out)
  );

  //Wire declarations for instance 'or_157' (Module coreir_or)
  wire [15:0] or_157__in0;
  wire [15:0] or_157__in1;
  wire [15:0] or_157__out;
  coreir_or #(.width(16)) or_157(
    .in0(or_157__in0),
    .in1(or_157__in1),
    .out(or_157__out)
  );

  //Wire declarations for instance 'or_159' (Module coreir_or)
  wire [15:0] or_159__in0;
  wire [15:0] or_159__in1;
  wire [15:0] or_159__out;
  coreir_or #(.width(16)) or_159(
    .in0(or_159__in0),
    .in1(or_159__in1),
    .out(or_159__out)
  );

  //Wire declarations for instance 'or_161' (Module coreir_or)
  wire [15:0] or_161__in0;
  wire [15:0] or_161__in1;
  wire [15:0] or_161__out;
  coreir_or #(.width(16)) or_161(
    .in0(or_161__in0),
    .in1(or_161__in1),
    .out(or_161__out)
  );

  //Wire declarations for instance 'or_163' (Module coreir_or)
  wire [15:0] or_163__in0;
  wire [15:0] or_163__in1;
  wire [15:0] or_163__out;
  coreir_or #(.width(16)) or_163(
    .in0(or_163__in0),
    .in1(or_163__in1),
    .out(or_163__out)
  );

  //Wire declarations for instance 'or_165' (Module coreir_or)
  wire [15:0] or_165__in0;
  wire [15:0] or_165__in1;
  wire [15:0] or_165__out;
  coreir_or #(.width(16)) or_165(
    .in0(or_165__in0),
    .in1(or_165__in1),
    .out(or_165__out)
  );

  //Wire declarations for instance 'or_167' (Module coreir_or)
  wire [15:0] or_167__in0;
  wire [15:0] or_167__in1;
  wire [15:0] or_167__out;
  coreir_or #(.width(16)) or_167(
    .in0(or_167__in0),
    .in1(or_167__in1),
    .out(or_167__out)
  );

  //Wire declarations for instance 'or_169' (Module coreir_or)
  wire [15:0] or_169__in0;
  wire [15:0] or_169__in1;
  wire [15:0] or_169__out;
  coreir_or #(.width(16)) or_169(
    .in0(or_169__in0),
    .in1(or_169__in1),
    .out(or_169__out)
  );

  //Wire declarations for instance 'or_17' (Module coreir_or)
  wire [15:0] or_17__in0;
  wire [15:0] or_17__in1;
  wire [15:0] or_17__out;
  coreir_or #(.width(16)) or_17(
    .in0(or_17__in0),
    .in1(or_17__in1),
    .out(or_17__out)
  );

  //Wire declarations for instance 'or_171' (Module coreir_or)
  wire [15:0] or_171__in0;
  wire [15:0] or_171__in1;
  wire [15:0] or_171__out;
  coreir_or #(.width(16)) or_171(
    .in0(or_171__in0),
    .in1(or_171__in1),
    .out(or_171__out)
  );

  //Wire declarations for instance 'or_173' (Module coreir_or)
  wire [15:0] or_173__in0;
  wire [15:0] or_173__in1;
  wire [15:0] or_173__out;
  coreir_or #(.width(16)) or_173(
    .in0(or_173__in0),
    .in1(or_173__in1),
    .out(or_173__out)
  );

  //Wire declarations for instance 'or_175' (Module coreir_or)
  wire [15:0] or_175__in0;
  wire [15:0] or_175__in1;
  wire [15:0] or_175__out;
  coreir_or #(.width(16)) or_175(
    .in0(or_175__in0),
    .in1(or_175__in1),
    .out(or_175__out)
  );

  //Wire declarations for instance 'or_177' (Module coreir_or)
  wire [15:0] or_177__in0;
  wire [15:0] or_177__in1;
  wire [15:0] or_177__out;
  coreir_or #(.width(16)) or_177(
    .in0(or_177__in0),
    .in1(or_177__in1),
    .out(or_177__out)
  );

  //Wire declarations for instance 'or_179' (Module coreir_or)
  wire [15:0] or_179__in0;
  wire [15:0] or_179__in1;
  wire [15:0] or_179__out;
  coreir_or #(.width(16)) or_179(
    .in0(or_179__in0),
    .in1(or_179__in1),
    .out(or_179__out)
  );

  //Wire declarations for instance 'or_181' (Module coreir_or)
  wire [15:0] or_181__in0;
  wire [15:0] or_181__in1;
  wire [15:0] or_181__out;
  coreir_or #(.width(16)) or_181(
    .in0(or_181__in0),
    .in1(or_181__in1),
    .out(or_181__out)
  );

  //Wire declarations for instance 'or_183' (Module coreir_or)
  wire [15:0] or_183__in0;
  wire [15:0] or_183__in1;
  wire [15:0] or_183__out;
  coreir_or #(.width(16)) or_183(
    .in0(or_183__in0),
    .in1(or_183__in1),
    .out(or_183__out)
  );

  //Wire declarations for instance 'or_185' (Module coreir_or)
  wire [15:0] or_185__in0;
  wire [15:0] or_185__in1;
  wire [15:0] or_185__out;
  coreir_or #(.width(16)) or_185(
    .in0(or_185__in0),
    .in1(or_185__in1),
    .out(or_185__out)
  );

  //Wire declarations for instance 'or_187' (Module coreir_or)
  wire [15:0] or_187__in0;
  wire [15:0] or_187__in1;
  wire [15:0] or_187__out;
  coreir_or #(.width(16)) or_187(
    .in0(or_187__in0),
    .in1(or_187__in1),
    .out(or_187__out)
  );

  //Wire declarations for instance 'or_189' (Module coreir_or)
  wire [15:0] or_189__in0;
  wire [15:0] or_189__in1;
  wire [15:0] or_189__out;
  coreir_or #(.width(16)) or_189(
    .in0(or_189__in0),
    .in1(or_189__in1),
    .out(or_189__out)
  );

  //Wire declarations for instance 'or_19' (Module coreir_or)
  wire [15:0] or_19__in0;
  wire [15:0] or_19__in1;
  wire [15:0] or_19__out;
  coreir_or #(.width(16)) or_19(
    .in0(or_19__in0),
    .in1(or_19__in1),
    .out(or_19__out)
  );

  //Wire declarations for instance 'or_191' (Module coreir_or)
  wire [15:0] or_191__in0;
  wire [15:0] or_191__in1;
  wire [15:0] or_191__out;
  coreir_or #(.width(16)) or_191(
    .in0(or_191__in0),
    .in1(or_191__in1),
    .out(or_191__out)
  );

  //Wire declarations for instance 'or_193' (Module coreir_or)
  wire [15:0] or_193__in0;
  wire [15:0] or_193__in1;
  wire [15:0] or_193__out;
  coreir_or #(.width(16)) or_193(
    .in0(or_193__in0),
    .in1(or_193__in1),
    .out(or_193__out)
  );

  //Wire declarations for instance 'or_195' (Module coreir_or)
  wire [15:0] or_195__in0;
  wire [15:0] or_195__in1;
  wire [15:0] or_195__out;
  coreir_or #(.width(16)) or_195(
    .in0(or_195__in0),
    .in1(or_195__in1),
    .out(or_195__out)
  );

  //Wire declarations for instance 'or_197' (Module coreir_or)
  wire [15:0] or_197__in0;
  wire [15:0] or_197__in1;
  wire [15:0] or_197__out;
  coreir_or #(.width(16)) or_197(
    .in0(or_197__in0),
    .in1(or_197__in1),
    .out(or_197__out)
  );

  //Wire declarations for instance 'or_199' (Module coreir_or)
  wire [15:0] or_199__in0;
  wire [15:0] or_199__in1;
  wire [15:0] or_199__out;
  coreir_or #(.width(16)) or_199(
    .in0(or_199__in0),
    .in1(or_199__in1),
    .out(or_199__out)
  );

  //Wire declarations for instance 'or_201' (Module coreir_or)
  wire [15:0] or_201__in0;
  wire [15:0] or_201__in1;
  wire [15:0] or_201__out;
  coreir_or #(.width(16)) or_201(
    .in0(or_201__in0),
    .in1(or_201__in1),
    .out(or_201__out)
  );

  //Wire declarations for instance 'or_203' (Module coreir_or)
  wire [15:0] or_203__in0;
  wire [15:0] or_203__in1;
  wire [15:0] or_203__out;
  coreir_or #(.width(16)) or_203(
    .in0(or_203__in0),
    .in1(or_203__in1),
    .out(or_203__out)
  );

  //Wire declarations for instance 'or_205' (Module coreir_or)
  wire [15:0] or_205__in0;
  wire [15:0] or_205__in1;
  wire [15:0] or_205__out;
  coreir_or #(.width(16)) or_205(
    .in0(or_205__in0),
    .in1(or_205__in1),
    .out(or_205__out)
  );

  //Wire declarations for instance 'or_207' (Module coreir_or)
  wire [15:0] or_207__in0;
  wire [15:0] or_207__in1;
  wire [15:0] or_207__out;
  coreir_or #(.width(16)) or_207(
    .in0(or_207__in0),
    .in1(or_207__in1),
    .out(or_207__out)
  );

  //Wire declarations for instance 'or_209' (Module coreir_or)
  wire [15:0] or_209__in0;
  wire [15:0] or_209__in1;
  wire [15:0] or_209__out;
  coreir_or #(.width(16)) or_209(
    .in0(or_209__in0),
    .in1(or_209__in1),
    .out(or_209__out)
  );

  //Wire declarations for instance 'or_21' (Module coreir_or)
  wire [15:0] or_21__in0;
  wire [15:0] or_21__in1;
  wire [15:0] or_21__out;
  coreir_or #(.width(16)) or_21(
    .in0(or_21__in0),
    .in1(or_21__in1),
    .out(or_21__out)
  );

  //Wire declarations for instance 'or_211' (Module coreir_or)
  wire [15:0] or_211__in0;
  wire [15:0] or_211__in1;
  wire [15:0] or_211__out;
  coreir_or #(.width(16)) or_211(
    .in0(or_211__in0),
    .in1(or_211__in1),
    .out(or_211__out)
  );

  //Wire declarations for instance 'or_213' (Module coreir_or)
  wire [15:0] or_213__in0;
  wire [15:0] or_213__in1;
  wire [15:0] or_213__out;
  coreir_or #(.width(16)) or_213(
    .in0(or_213__in0),
    .in1(or_213__in1),
    .out(or_213__out)
  );

  //Wire declarations for instance 'or_215' (Module coreir_or)
  wire [15:0] or_215__in0;
  wire [15:0] or_215__in1;
  wire [15:0] or_215__out;
  coreir_or #(.width(16)) or_215(
    .in0(or_215__in0),
    .in1(or_215__in1),
    .out(or_215__out)
  );

  //Wire declarations for instance 'or_217' (Module coreir_or)
  wire [15:0] or_217__in0;
  wire [15:0] or_217__in1;
  wire [15:0] or_217__out;
  coreir_or #(.width(16)) or_217(
    .in0(or_217__in0),
    .in1(or_217__in1),
    .out(or_217__out)
  );

  //Wire declarations for instance 'or_219' (Module coreir_or)
  wire [15:0] or_219__in0;
  wire [15:0] or_219__in1;
  wire [15:0] or_219__out;
  coreir_or #(.width(16)) or_219(
    .in0(or_219__in0),
    .in1(or_219__in1),
    .out(or_219__out)
  );

  //Wire declarations for instance 'or_221' (Module coreir_or)
  wire [15:0] or_221__in0;
  wire [15:0] or_221__in1;
  wire [15:0] or_221__out;
  coreir_or #(.width(16)) or_221(
    .in0(or_221__in0),
    .in1(or_221__in1),
    .out(or_221__out)
  );

  //Wire declarations for instance 'or_223' (Module coreir_or)
  wire [15:0] or_223__in0;
  wire [15:0] or_223__in1;
  wire [15:0] or_223__out;
  coreir_or #(.width(16)) or_223(
    .in0(or_223__in0),
    .in1(or_223__in1),
    .out(or_223__out)
  );

  //Wire declarations for instance 'or_225' (Module coreir_or)
  wire [15:0] or_225__in0;
  wire [15:0] or_225__in1;
  wire [15:0] or_225__out;
  coreir_or #(.width(16)) or_225(
    .in0(or_225__in0),
    .in1(or_225__in1),
    .out(or_225__out)
  );

  //Wire declarations for instance 'or_227' (Module coreir_or)
  wire [15:0] or_227__in0;
  wire [15:0] or_227__in1;
  wire [15:0] or_227__out;
  coreir_or #(.width(16)) or_227(
    .in0(or_227__in0),
    .in1(or_227__in1),
    .out(or_227__out)
  );

  //Wire declarations for instance 'or_229' (Module coreir_or)
  wire [15:0] or_229__in0;
  wire [15:0] or_229__in1;
  wire [15:0] or_229__out;
  coreir_or #(.width(16)) or_229(
    .in0(or_229__in0),
    .in1(or_229__in1),
    .out(or_229__out)
  );

  //Wire declarations for instance 'or_23' (Module coreir_or)
  wire [15:0] or_23__in0;
  wire [15:0] or_23__in1;
  wire [15:0] or_23__out;
  coreir_or #(.width(16)) or_23(
    .in0(or_23__in0),
    .in1(or_23__in1),
    .out(or_23__out)
  );

  //Wire declarations for instance 'or_231' (Module coreir_or)
  wire [15:0] or_231__in0;
  wire [15:0] or_231__in1;
  wire [15:0] or_231__out;
  coreir_or #(.width(16)) or_231(
    .in0(or_231__in0),
    .in1(or_231__in1),
    .out(or_231__out)
  );

  //Wire declarations for instance 'or_233' (Module coreir_or)
  wire [15:0] or_233__in0;
  wire [15:0] or_233__in1;
  wire [15:0] or_233__out;
  coreir_or #(.width(16)) or_233(
    .in0(or_233__in0),
    .in1(or_233__in1),
    .out(or_233__out)
  );

  //Wire declarations for instance 'or_235' (Module coreir_or)
  wire [15:0] or_235__in0;
  wire [15:0] or_235__in1;
  wire [15:0] or_235__out;
  coreir_or #(.width(16)) or_235(
    .in0(or_235__in0),
    .in1(or_235__in1),
    .out(or_235__out)
  );

  //Wire declarations for instance 'or_237' (Module coreir_or)
  wire [15:0] or_237__in0;
  wire [15:0] or_237__in1;
  wire [15:0] or_237__out;
  coreir_or #(.width(16)) or_237(
    .in0(or_237__in0),
    .in1(or_237__in1),
    .out(or_237__out)
  );

  //Wire declarations for instance 'or_239' (Module coreir_or)
  wire [15:0] or_239__in0;
  wire [15:0] or_239__in1;
  wire [15:0] or_239__out;
  coreir_or #(.width(16)) or_239(
    .in0(or_239__in0),
    .in1(or_239__in1),
    .out(or_239__out)
  );

  //Wire declarations for instance 'or_241' (Module coreir_or)
  wire [15:0] or_241__in0;
  wire [15:0] or_241__in1;
  wire [15:0] or_241__out;
  coreir_or #(.width(16)) or_241(
    .in0(or_241__in0),
    .in1(or_241__in1),
    .out(or_241__out)
  );

  //Wire declarations for instance 'or_243' (Module coreir_or)
  wire [15:0] or_243__in0;
  wire [15:0] or_243__in1;
  wire [15:0] or_243__out;
  coreir_or #(.width(16)) or_243(
    .in0(or_243__in0),
    .in1(or_243__in1),
    .out(or_243__out)
  );

  //Wire declarations for instance 'or_245' (Module coreir_or)
  wire [15:0] or_245__in0;
  wire [15:0] or_245__in1;
  wire [15:0] or_245__out;
  coreir_or #(.width(16)) or_245(
    .in0(or_245__in0),
    .in1(or_245__in1),
    .out(or_245__out)
  );

  //Wire declarations for instance 'or_247' (Module coreir_or)
  wire [15:0] or_247__in0;
  wire [15:0] or_247__in1;
  wire [15:0] or_247__out;
  coreir_or #(.width(16)) or_247(
    .in0(or_247__in0),
    .in1(or_247__in1),
    .out(or_247__out)
  );

  //Wire declarations for instance 'or_249' (Module coreir_or)
  wire [15:0] or_249__in0;
  wire [15:0] or_249__in1;
  wire [15:0] or_249__out;
  coreir_or #(.width(16)) or_249(
    .in0(or_249__in0),
    .in1(or_249__in1),
    .out(or_249__out)
  );

  //Wire declarations for instance 'or_25' (Module coreir_or)
  wire [15:0] or_25__in0;
  wire [15:0] or_25__in1;
  wire [15:0] or_25__out;
  coreir_or #(.width(16)) or_25(
    .in0(or_25__in0),
    .in1(or_25__in1),
    .out(or_25__out)
  );

  //Wire declarations for instance 'or_251' (Module coreir_or)
  wire [15:0] or_251__in0;
  wire [15:0] or_251__in1;
  wire [15:0] or_251__out;
  coreir_or #(.width(16)) or_251(
    .in0(or_251__in0),
    .in1(or_251__in1),
    .out(or_251__out)
  );

  //Wire declarations for instance 'or_253' (Module coreir_or)
  wire [15:0] or_253__in0;
  wire [15:0] or_253__in1;
  wire [15:0] or_253__out;
  coreir_or #(.width(16)) or_253(
    .in0(or_253__in0),
    .in1(or_253__in1),
    .out(or_253__out)
  );

  //Wire declarations for instance 'or_255' (Module coreir_or)
  wire [15:0] or_255__in0;
  wire [15:0] or_255__in1;
  wire [15:0] or_255__out;
  coreir_or #(.width(16)) or_255(
    .in0(or_255__in0),
    .in1(or_255__in1),
    .out(or_255__out)
  );

  //Wire declarations for instance 'or_257' (Module coreir_or)
  wire [15:0] or_257__in0;
  wire [15:0] or_257__in1;
  wire [15:0] or_257__out;
  coreir_or #(.width(16)) or_257(
    .in0(or_257__in0),
    .in1(or_257__in1),
    .out(or_257__out)
  );

  //Wire declarations for instance 'or_259' (Module coreir_or)
  wire [15:0] or_259__in0;
  wire [15:0] or_259__in1;
  wire [15:0] or_259__out;
  coreir_or #(.width(16)) or_259(
    .in0(or_259__in0),
    .in1(or_259__in1),
    .out(or_259__out)
  );

  //Wire declarations for instance 'or_261' (Module coreir_or)
  wire [15:0] or_261__in0;
  wire [15:0] or_261__in1;
  wire [15:0] or_261__out;
  coreir_or #(.width(16)) or_261(
    .in0(or_261__in0),
    .in1(or_261__in1),
    .out(or_261__out)
  );

  //Wire declarations for instance 'or_263' (Module coreir_or)
  wire [15:0] or_263__in0;
  wire [15:0] or_263__in1;
  wire [15:0] or_263__out;
  coreir_or #(.width(16)) or_263(
    .in0(or_263__in0),
    .in1(or_263__in1),
    .out(or_263__out)
  );

  //Wire declarations for instance 'or_265' (Module coreir_or)
  wire [15:0] or_265__in0;
  wire [15:0] or_265__in1;
  wire [15:0] or_265__out;
  coreir_or #(.width(16)) or_265(
    .in0(or_265__in0),
    .in1(or_265__in1),
    .out(or_265__out)
  );

  //Wire declarations for instance 'or_267' (Module coreir_or)
  wire [15:0] or_267__in0;
  wire [15:0] or_267__in1;
  wire [15:0] or_267__out;
  coreir_or #(.width(16)) or_267(
    .in0(or_267__in0),
    .in1(or_267__in1),
    .out(or_267__out)
  );

  //Wire declarations for instance 'or_269' (Module coreir_or)
  wire [15:0] or_269__in0;
  wire [15:0] or_269__in1;
  wire [15:0] or_269__out;
  coreir_or #(.width(16)) or_269(
    .in0(or_269__in0),
    .in1(or_269__in1),
    .out(or_269__out)
  );

  //Wire declarations for instance 'or_27' (Module coreir_or)
  wire [15:0] or_27__in0;
  wire [15:0] or_27__in1;
  wire [15:0] or_27__out;
  coreir_or #(.width(16)) or_27(
    .in0(or_27__in0),
    .in1(or_27__in1),
    .out(or_27__out)
  );

  //Wire declarations for instance 'or_271' (Module coreir_or)
  wire [15:0] or_271__in0;
  wire [15:0] or_271__in1;
  wire [15:0] or_271__out;
  coreir_or #(.width(16)) or_271(
    .in0(or_271__in0),
    .in1(or_271__in1),
    .out(or_271__out)
  );

  //Wire declarations for instance 'or_273' (Module coreir_or)
  wire [15:0] or_273__in0;
  wire [15:0] or_273__in1;
  wire [15:0] or_273__out;
  coreir_or #(.width(16)) or_273(
    .in0(or_273__in0),
    .in1(or_273__in1),
    .out(or_273__out)
  );

  //Wire declarations for instance 'or_275' (Module coreir_or)
  wire [15:0] or_275__in0;
  wire [15:0] or_275__in1;
  wire [15:0] or_275__out;
  coreir_or #(.width(16)) or_275(
    .in0(or_275__in0),
    .in1(or_275__in1),
    .out(or_275__out)
  );

  //Wire declarations for instance 'or_277' (Module coreir_or)
  wire [15:0] or_277__in0;
  wire [15:0] or_277__in1;
  wire [15:0] or_277__out;
  coreir_or #(.width(16)) or_277(
    .in0(or_277__in0),
    .in1(or_277__in1),
    .out(or_277__out)
  );

  //Wire declarations for instance 'or_279' (Module coreir_or)
  wire [15:0] or_279__in0;
  wire [15:0] or_279__in1;
  wire [15:0] or_279__out;
  coreir_or #(.width(16)) or_279(
    .in0(or_279__in0),
    .in1(or_279__in1),
    .out(or_279__out)
  );

  //Wire declarations for instance 'or_281' (Module coreir_or)
  wire [15:0] or_281__in0;
  wire [15:0] or_281__in1;
  wire [15:0] or_281__out;
  coreir_or #(.width(16)) or_281(
    .in0(or_281__in0),
    .in1(or_281__in1),
    .out(or_281__out)
  );

  //Wire declarations for instance 'or_283' (Module coreir_or)
  wire [15:0] or_283__in0;
  wire [15:0] or_283__in1;
  wire [15:0] or_283__out;
  coreir_or #(.width(16)) or_283(
    .in0(or_283__in0),
    .in1(or_283__in1),
    .out(or_283__out)
  );

  //Wire declarations for instance 'or_285' (Module coreir_or)
  wire [15:0] or_285__in0;
  wire [15:0] or_285__in1;
  wire [15:0] or_285__out;
  coreir_or #(.width(16)) or_285(
    .in0(or_285__in0),
    .in1(or_285__in1),
    .out(or_285__out)
  );

  //Wire declarations for instance 'or_287' (Module coreir_or)
  wire [15:0] or_287__in0;
  wire [15:0] or_287__in1;
  wire [15:0] or_287__out;
  coreir_or #(.width(16)) or_287(
    .in0(or_287__in0),
    .in1(or_287__in1),
    .out(or_287__out)
  );

  //Wire declarations for instance 'or_289' (Module coreir_or)
  wire [15:0] or_289__in0;
  wire [15:0] or_289__in1;
  wire [15:0] or_289__out;
  coreir_or #(.width(16)) or_289(
    .in0(or_289__in0),
    .in1(or_289__in1),
    .out(or_289__out)
  );

  //Wire declarations for instance 'or_29' (Module coreir_or)
  wire [15:0] or_29__in0;
  wire [15:0] or_29__in1;
  wire [15:0] or_29__out;
  coreir_or #(.width(16)) or_29(
    .in0(or_29__in0),
    .in1(or_29__in1),
    .out(or_29__out)
  );

  //Wire declarations for instance 'or_291' (Module coreir_or)
  wire [15:0] or_291__in0;
  wire [15:0] or_291__in1;
  wire [15:0] or_291__out;
  coreir_or #(.width(16)) or_291(
    .in0(or_291__in0),
    .in1(or_291__in1),
    .out(or_291__out)
  );

  //Wire declarations for instance 'or_293' (Module coreir_or)
  wire [15:0] or_293__in0;
  wire [15:0] or_293__in1;
  wire [15:0] or_293__out;
  coreir_or #(.width(16)) or_293(
    .in0(or_293__in0),
    .in1(or_293__in1),
    .out(or_293__out)
  );

  //Wire declarations for instance 'or_295' (Module coreir_or)
  wire [15:0] or_295__in0;
  wire [15:0] or_295__in1;
  wire [15:0] or_295__out;
  coreir_or #(.width(16)) or_295(
    .in0(or_295__in0),
    .in1(or_295__in1),
    .out(or_295__out)
  );

  //Wire declarations for instance 'or_297' (Module coreir_or)
  wire [15:0] or_297__in0;
  wire [15:0] or_297__in1;
  wire [15:0] or_297__out;
  coreir_or #(.width(16)) or_297(
    .in0(or_297__in0),
    .in1(or_297__in1),
    .out(or_297__out)
  );

  //Wire declarations for instance 'or_299' (Module coreir_or)
  wire [15:0] or_299__in0;
  wire [15:0] or_299__in1;
  wire [15:0] or_299__out;
  coreir_or #(.width(16)) or_299(
    .in0(or_299__in0),
    .in1(or_299__in1),
    .out(or_299__out)
  );

  //Wire declarations for instance 'or_3' (Module coreir_or)
  wire [15:0] or_3__in0;
  wire [15:0] or_3__in1;
  wire [15:0] or_3__out;
  coreir_or #(.width(16)) or_3(
    .in0(or_3__in0),
    .in1(or_3__in1),
    .out(or_3__out)
  );

  //Wire declarations for instance 'or_301' (Module coreir_or)
  wire [15:0] or_301__in0;
  wire [15:0] or_301__in1;
  wire [15:0] or_301__out;
  coreir_or #(.width(16)) or_301(
    .in0(or_301__in0),
    .in1(or_301__in1),
    .out(or_301__out)
  );

  //Wire declarations for instance 'or_303' (Module coreir_or)
  wire [15:0] or_303__in0;
  wire [15:0] or_303__in1;
  wire [15:0] or_303__out;
  coreir_or #(.width(16)) or_303(
    .in0(or_303__in0),
    .in1(or_303__in1),
    .out(or_303__out)
  );

  //Wire declarations for instance 'or_305' (Module coreir_or)
  wire [15:0] or_305__in0;
  wire [15:0] or_305__in1;
  wire [15:0] or_305__out;
  coreir_or #(.width(16)) or_305(
    .in0(or_305__in0),
    .in1(or_305__in1),
    .out(or_305__out)
  );

  //Wire declarations for instance 'or_307' (Module coreir_or)
  wire [15:0] or_307__in0;
  wire [15:0] or_307__in1;
  wire [15:0] or_307__out;
  coreir_or #(.width(16)) or_307(
    .in0(or_307__in0),
    .in1(or_307__in1),
    .out(or_307__out)
  );

  //Wire declarations for instance 'or_309' (Module coreir_or)
  wire [15:0] or_309__in0;
  wire [15:0] or_309__in1;
  wire [15:0] or_309__out;
  coreir_or #(.width(16)) or_309(
    .in0(or_309__in0),
    .in1(or_309__in1),
    .out(or_309__out)
  );

  //Wire declarations for instance 'or_31' (Module coreir_or)
  wire [15:0] or_31__in0;
  wire [15:0] or_31__in1;
  wire [15:0] or_31__out;
  coreir_or #(.width(16)) or_31(
    .in0(or_31__in0),
    .in1(or_31__in1),
    .out(or_31__out)
  );

  //Wire declarations for instance 'or_311' (Module coreir_or)
  wire [15:0] or_311__in0;
  wire [15:0] or_311__in1;
  wire [15:0] or_311__out;
  coreir_or #(.width(16)) or_311(
    .in0(or_311__in0),
    .in1(or_311__in1),
    .out(or_311__out)
  );

  //Wire declarations for instance 'or_313' (Module coreir_or)
  wire [15:0] or_313__in0;
  wire [15:0] or_313__in1;
  wire [15:0] or_313__out;
  coreir_or #(.width(16)) or_313(
    .in0(or_313__in0),
    .in1(or_313__in1),
    .out(or_313__out)
  );

  //Wire declarations for instance 'or_315' (Module coreir_or)
  wire [15:0] or_315__in0;
  wire [15:0] or_315__in1;
  wire [15:0] or_315__out;
  coreir_or #(.width(16)) or_315(
    .in0(or_315__in0),
    .in1(or_315__in1),
    .out(or_315__out)
  );

  //Wire declarations for instance 'or_317' (Module coreir_or)
  wire [15:0] or_317__in0;
  wire [15:0] or_317__in1;
  wire [15:0] or_317__out;
  coreir_or #(.width(16)) or_317(
    .in0(or_317__in0),
    .in1(or_317__in1),
    .out(or_317__out)
  );

  //Wire declarations for instance 'or_319' (Module coreir_or)
  wire [15:0] or_319__in0;
  wire [15:0] or_319__in1;
  wire [15:0] or_319__out;
  coreir_or #(.width(16)) or_319(
    .in0(or_319__in0),
    .in1(or_319__in1),
    .out(or_319__out)
  );

  //Wire declarations for instance 'or_321' (Module coreir_or)
  wire [15:0] or_321__in0;
  wire [15:0] or_321__in1;
  wire [15:0] or_321__out;
  coreir_or #(.width(16)) or_321(
    .in0(or_321__in0),
    .in1(or_321__in1),
    .out(or_321__out)
  );

  //Wire declarations for instance 'or_323' (Module coreir_or)
  wire [15:0] or_323__in0;
  wire [15:0] or_323__in1;
  wire [15:0] or_323__out;
  coreir_or #(.width(16)) or_323(
    .in0(or_323__in0),
    .in1(or_323__in1),
    .out(or_323__out)
  );

  //Wire declarations for instance 'or_325' (Module coreir_or)
  wire [15:0] or_325__in0;
  wire [15:0] or_325__in1;
  wire [15:0] or_325__out;
  coreir_or #(.width(16)) or_325(
    .in0(or_325__in0),
    .in1(or_325__in1),
    .out(or_325__out)
  );

  //Wire declarations for instance 'or_327' (Module coreir_or)
  wire [15:0] or_327__in0;
  wire [15:0] or_327__in1;
  wire [15:0] or_327__out;
  coreir_or #(.width(16)) or_327(
    .in0(or_327__in0),
    .in1(or_327__in1),
    .out(or_327__out)
  );

  //Wire declarations for instance 'or_329' (Module coreir_or)
  wire [15:0] or_329__in0;
  wire [15:0] or_329__in1;
  wire [15:0] or_329__out;
  coreir_or #(.width(16)) or_329(
    .in0(or_329__in0),
    .in1(or_329__in1),
    .out(or_329__out)
  );

  //Wire declarations for instance 'or_33' (Module coreir_or)
  wire [15:0] or_33__in0;
  wire [15:0] or_33__in1;
  wire [15:0] or_33__out;
  coreir_or #(.width(16)) or_33(
    .in0(or_33__in0),
    .in1(or_33__in1),
    .out(or_33__out)
  );

  //Wire declarations for instance 'or_331' (Module coreir_or)
  wire [15:0] or_331__in0;
  wire [15:0] or_331__in1;
  wire [15:0] or_331__out;
  coreir_or #(.width(16)) or_331(
    .in0(or_331__in0),
    .in1(or_331__in1),
    .out(or_331__out)
  );

  //Wire declarations for instance 'or_333' (Module coreir_or)
  wire [15:0] or_333__in0;
  wire [15:0] or_333__in1;
  wire [15:0] or_333__out;
  coreir_or #(.width(16)) or_333(
    .in0(or_333__in0),
    .in1(or_333__in1),
    .out(or_333__out)
  );

  //Wire declarations for instance 'or_335' (Module coreir_or)
  wire [15:0] or_335__in0;
  wire [15:0] or_335__in1;
  wire [15:0] or_335__out;
  coreir_or #(.width(16)) or_335(
    .in0(or_335__in0),
    .in1(or_335__in1),
    .out(or_335__out)
  );

  //Wire declarations for instance 'or_337' (Module coreir_or)
  wire [15:0] or_337__in0;
  wire [15:0] or_337__in1;
  wire [15:0] or_337__out;
  coreir_or #(.width(16)) or_337(
    .in0(or_337__in0),
    .in1(or_337__in1),
    .out(or_337__out)
  );

  //Wire declarations for instance 'or_339' (Module coreir_or)
  wire [15:0] or_339__in0;
  wire [15:0] or_339__in1;
  wire [15:0] or_339__out;
  coreir_or #(.width(16)) or_339(
    .in0(or_339__in0),
    .in1(or_339__in1),
    .out(or_339__out)
  );

  //Wire declarations for instance 'or_341' (Module coreir_or)
  wire [15:0] or_341__in0;
  wire [15:0] or_341__in1;
  wire [15:0] or_341__out;
  coreir_or #(.width(16)) or_341(
    .in0(or_341__in0),
    .in1(or_341__in1),
    .out(or_341__out)
  );

  //Wire declarations for instance 'or_343' (Module coreir_or)
  wire [15:0] or_343__in0;
  wire [15:0] or_343__in1;
  wire [15:0] or_343__out;
  coreir_or #(.width(16)) or_343(
    .in0(or_343__in0),
    .in1(or_343__in1),
    .out(or_343__out)
  );

  //Wire declarations for instance 'or_345' (Module coreir_or)
  wire [15:0] or_345__in0;
  wire [15:0] or_345__in1;
  wire [15:0] or_345__out;
  coreir_or #(.width(16)) or_345(
    .in0(or_345__in0),
    .in1(or_345__in1),
    .out(or_345__out)
  );

  //Wire declarations for instance 'or_347' (Module coreir_or)
  wire [15:0] or_347__in0;
  wire [15:0] or_347__in1;
  wire [15:0] or_347__out;
  coreir_or #(.width(16)) or_347(
    .in0(or_347__in0),
    .in1(or_347__in1),
    .out(or_347__out)
  );

  //Wire declarations for instance 'or_349' (Module coreir_or)
  wire [15:0] or_349__in0;
  wire [15:0] or_349__in1;
  wire [15:0] or_349__out;
  coreir_or #(.width(16)) or_349(
    .in0(or_349__in0),
    .in1(or_349__in1),
    .out(or_349__out)
  );

  //Wire declarations for instance 'or_35' (Module coreir_or)
  wire [15:0] or_35__in0;
  wire [15:0] or_35__in1;
  wire [15:0] or_35__out;
  coreir_or #(.width(16)) or_35(
    .in0(or_35__in0),
    .in1(or_35__in1),
    .out(or_35__out)
  );

  //Wire declarations for instance 'or_351' (Module coreir_or)
  wire [15:0] or_351__in0;
  wire [15:0] or_351__in1;
  wire [15:0] or_351__out;
  coreir_or #(.width(16)) or_351(
    .in0(or_351__in0),
    .in1(or_351__in1),
    .out(or_351__out)
  );

  //Wire declarations for instance 'or_353' (Module coreir_or)
  wire [15:0] or_353__in0;
  wire [15:0] or_353__in1;
  wire [15:0] or_353__out;
  coreir_or #(.width(16)) or_353(
    .in0(or_353__in0),
    .in1(or_353__in1),
    .out(or_353__out)
  );

  //Wire declarations for instance 'or_355' (Module coreir_or)
  wire [15:0] or_355__in0;
  wire [15:0] or_355__in1;
  wire [15:0] or_355__out;
  coreir_or #(.width(16)) or_355(
    .in0(or_355__in0),
    .in1(or_355__in1),
    .out(or_355__out)
  );

  //Wire declarations for instance 'or_357' (Module coreir_or)
  wire [15:0] or_357__in0;
  wire [15:0] or_357__in1;
  wire [15:0] or_357__out;
  coreir_or #(.width(16)) or_357(
    .in0(or_357__in0),
    .in1(or_357__in1),
    .out(or_357__out)
  );

  //Wire declarations for instance 'or_359' (Module coreir_or)
  wire [15:0] or_359__in0;
  wire [15:0] or_359__in1;
  wire [15:0] or_359__out;
  coreir_or #(.width(16)) or_359(
    .in0(or_359__in0),
    .in1(or_359__in1),
    .out(or_359__out)
  );

  //Wire declarations for instance 'or_361' (Module coreir_or)
  wire [15:0] or_361__in0;
  wire [15:0] or_361__in1;
  wire [15:0] or_361__out;
  coreir_or #(.width(16)) or_361(
    .in0(or_361__in0),
    .in1(or_361__in1),
    .out(or_361__out)
  );

  //Wire declarations for instance 'or_363' (Module coreir_or)
  wire [15:0] or_363__in0;
  wire [15:0] or_363__in1;
  wire [15:0] or_363__out;
  coreir_or #(.width(16)) or_363(
    .in0(or_363__in0),
    .in1(or_363__in1),
    .out(or_363__out)
  );

  //Wire declarations for instance 'or_365' (Module coreir_or)
  wire [15:0] or_365__in0;
  wire [15:0] or_365__in1;
  wire [15:0] or_365__out;
  coreir_or #(.width(16)) or_365(
    .in0(or_365__in0),
    .in1(or_365__in1),
    .out(or_365__out)
  );

  //Wire declarations for instance 'or_367' (Module coreir_or)
  wire [15:0] or_367__in0;
  wire [15:0] or_367__in1;
  wire [15:0] or_367__out;
  coreir_or #(.width(16)) or_367(
    .in0(or_367__in0),
    .in1(or_367__in1),
    .out(or_367__out)
  );

  //Wire declarations for instance 'or_369' (Module coreir_or)
  wire [15:0] or_369__in0;
  wire [15:0] or_369__in1;
  wire [15:0] or_369__out;
  coreir_or #(.width(16)) or_369(
    .in0(or_369__in0),
    .in1(or_369__in1),
    .out(or_369__out)
  );

  //Wire declarations for instance 'or_37' (Module coreir_or)
  wire [15:0] or_37__in0;
  wire [15:0] or_37__in1;
  wire [15:0] or_37__out;
  coreir_or #(.width(16)) or_37(
    .in0(or_37__in0),
    .in1(or_37__in1),
    .out(or_37__out)
  );

  //Wire declarations for instance 'or_371' (Module coreir_or)
  wire [15:0] or_371__in0;
  wire [15:0] or_371__in1;
  wire [15:0] or_371__out;
  coreir_or #(.width(16)) or_371(
    .in0(or_371__in0),
    .in1(or_371__in1),
    .out(or_371__out)
  );

  //Wire declarations for instance 'or_373' (Module coreir_or)
  wire [15:0] or_373__in0;
  wire [15:0] or_373__in1;
  wire [15:0] or_373__out;
  coreir_or #(.width(16)) or_373(
    .in0(or_373__in0),
    .in1(or_373__in1),
    .out(or_373__out)
  );

  //Wire declarations for instance 'or_375' (Module coreir_or)
  wire [15:0] or_375__in0;
  wire [15:0] or_375__in1;
  wire [15:0] or_375__out;
  coreir_or #(.width(16)) or_375(
    .in0(or_375__in0),
    .in1(or_375__in1),
    .out(or_375__out)
  );

  //Wire declarations for instance 'or_377' (Module coreir_or)
  wire [15:0] or_377__in0;
  wire [15:0] or_377__in1;
  wire [15:0] or_377__out;
  coreir_or #(.width(16)) or_377(
    .in0(or_377__in0),
    .in1(or_377__in1),
    .out(or_377__out)
  );

  //Wire declarations for instance 'or_379' (Module coreir_or)
  wire [15:0] or_379__in0;
  wire [15:0] or_379__in1;
  wire [15:0] or_379__out;
  coreir_or #(.width(16)) or_379(
    .in0(or_379__in0),
    .in1(or_379__in1),
    .out(or_379__out)
  );

  //Wire declarations for instance 'or_381' (Module coreir_or)
  wire [15:0] or_381__in0;
  wire [15:0] or_381__in1;
  wire [15:0] or_381__out;
  coreir_or #(.width(16)) or_381(
    .in0(or_381__in0),
    .in1(or_381__in1),
    .out(or_381__out)
  );

  //Wire declarations for instance 'or_383' (Module coreir_or)
  wire [15:0] or_383__in0;
  wire [15:0] or_383__in1;
  wire [15:0] or_383__out;
  coreir_or #(.width(16)) or_383(
    .in0(or_383__in0),
    .in1(or_383__in1),
    .out(or_383__out)
  );

  //Wire declarations for instance 'or_385' (Module coreir_or)
  wire [15:0] or_385__in0;
  wire [15:0] or_385__in1;
  wire [15:0] or_385__out;
  coreir_or #(.width(16)) or_385(
    .in0(or_385__in0),
    .in1(or_385__in1),
    .out(or_385__out)
  );

  //Wire declarations for instance 'or_387' (Module coreir_or)
  wire [15:0] or_387__in0;
  wire [15:0] or_387__in1;
  wire [15:0] or_387__out;
  coreir_or #(.width(16)) or_387(
    .in0(or_387__in0),
    .in1(or_387__in1),
    .out(or_387__out)
  );

  //Wire declarations for instance 'or_389' (Module coreir_or)
  wire [15:0] or_389__in0;
  wire [15:0] or_389__in1;
  wire [15:0] or_389__out;
  coreir_or #(.width(16)) or_389(
    .in0(or_389__in0),
    .in1(or_389__in1),
    .out(or_389__out)
  );

  //Wire declarations for instance 'or_39' (Module coreir_or)
  wire [15:0] or_39__in0;
  wire [15:0] or_39__in1;
  wire [15:0] or_39__out;
  coreir_or #(.width(16)) or_39(
    .in0(or_39__in0),
    .in1(or_39__in1),
    .out(or_39__out)
  );

  //Wire declarations for instance 'or_391' (Module coreir_or)
  wire [15:0] or_391__in0;
  wire [15:0] or_391__in1;
  wire [15:0] or_391__out;
  coreir_or #(.width(16)) or_391(
    .in0(or_391__in0),
    .in1(or_391__in1),
    .out(or_391__out)
  );

  //Wire declarations for instance 'or_393' (Module coreir_or)
  wire [15:0] or_393__in0;
  wire [15:0] or_393__in1;
  wire [15:0] or_393__out;
  coreir_or #(.width(16)) or_393(
    .in0(or_393__in0),
    .in1(or_393__in1),
    .out(or_393__out)
  );

  //Wire declarations for instance 'or_395' (Module coreir_or)
  wire [15:0] or_395__in0;
  wire [15:0] or_395__in1;
  wire [15:0] or_395__out;
  coreir_or #(.width(16)) or_395(
    .in0(or_395__in0),
    .in1(or_395__in1),
    .out(or_395__out)
  );

  //Wire declarations for instance 'or_397' (Module coreir_or)
  wire [15:0] or_397__in0;
  wire [15:0] or_397__in1;
  wire [15:0] or_397__out;
  coreir_or #(.width(16)) or_397(
    .in0(or_397__in0),
    .in1(or_397__in1),
    .out(or_397__out)
  );

  //Wire declarations for instance 'or_399' (Module coreir_or)
  wire [15:0] or_399__in0;
  wire [15:0] or_399__in1;
  wire [15:0] or_399__out;
  coreir_or #(.width(16)) or_399(
    .in0(or_399__in0),
    .in1(or_399__in1),
    .out(or_399__out)
  );

  //Wire declarations for instance 'or_401' (Module coreir_or)
  wire [15:0] or_401__in0;
  wire [15:0] or_401__in1;
  wire [15:0] or_401__out;
  coreir_or #(.width(16)) or_401(
    .in0(or_401__in0),
    .in1(or_401__in1),
    .out(or_401__out)
  );

  //Wire declarations for instance 'or_403' (Module coreir_or)
  wire [15:0] or_403__in0;
  wire [15:0] or_403__in1;
  wire [15:0] or_403__out;
  coreir_or #(.width(16)) or_403(
    .in0(or_403__in0),
    .in1(or_403__in1),
    .out(or_403__out)
  );

  //Wire declarations for instance 'or_405' (Module coreir_or)
  wire [15:0] or_405__in0;
  wire [15:0] or_405__in1;
  wire [15:0] or_405__out;
  coreir_or #(.width(16)) or_405(
    .in0(or_405__in0),
    .in1(or_405__in1),
    .out(or_405__out)
  );

  //Wire declarations for instance 'or_407' (Module coreir_or)
  wire [15:0] or_407__in0;
  wire [15:0] or_407__in1;
  wire [15:0] or_407__out;
  coreir_or #(.width(16)) or_407(
    .in0(or_407__in0),
    .in1(or_407__in1),
    .out(or_407__out)
  );

  //Wire declarations for instance 'or_409' (Module coreir_or)
  wire [15:0] or_409__in0;
  wire [15:0] or_409__in1;
  wire [15:0] or_409__out;
  coreir_or #(.width(16)) or_409(
    .in0(or_409__in0),
    .in1(or_409__in1),
    .out(or_409__out)
  );

  //Wire declarations for instance 'or_41' (Module coreir_or)
  wire [15:0] or_41__in0;
  wire [15:0] or_41__in1;
  wire [15:0] or_41__out;
  coreir_or #(.width(16)) or_41(
    .in0(or_41__in0),
    .in1(or_41__in1),
    .out(or_41__out)
  );

  //Wire declarations for instance 'or_411' (Module coreir_or)
  wire [15:0] or_411__in0;
  wire [15:0] or_411__in1;
  wire [15:0] or_411__out;
  coreir_or #(.width(16)) or_411(
    .in0(or_411__in0),
    .in1(or_411__in1),
    .out(or_411__out)
  );

  //Wire declarations for instance 'or_413' (Module coreir_or)
  wire [15:0] or_413__in0;
  wire [15:0] or_413__in1;
  wire [15:0] or_413__out;
  coreir_or #(.width(16)) or_413(
    .in0(or_413__in0),
    .in1(or_413__in1),
    .out(or_413__out)
  );

  //Wire declarations for instance 'or_415' (Module coreir_or)
  wire [15:0] or_415__in0;
  wire [15:0] or_415__in1;
  wire [15:0] or_415__out;
  coreir_or #(.width(16)) or_415(
    .in0(or_415__in0),
    .in1(or_415__in1),
    .out(or_415__out)
  );

  //Wire declarations for instance 'or_417' (Module coreir_or)
  wire [15:0] or_417__in0;
  wire [15:0] or_417__in1;
  wire [15:0] or_417__out;
  coreir_or #(.width(16)) or_417(
    .in0(or_417__in0),
    .in1(or_417__in1),
    .out(or_417__out)
  );

  //Wire declarations for instance 'or_419' (Module coreir_or)
  wire [15:0] or_419__in0;
  wire [15:0] or_419__in1;
  wire [15:0] or_419__out;
  coreir_or #(.width(16)) or_419(
    .in0(or_419__in0),
    .in1(or_419__in1),
    .out(or_419__out)
  );

  //Wire declarations for instance 'or_421' (Module coreir_or)
  wire [15:0] or_421__in0;
  wire [15:0] or_421__in1;
  wire [15:0] or_421__out;
  coreir_or #(.width(16)) or_421(
    .in0(or_421__in0),
    .in1(or_421__in1),
    .out(or_421__out)
  );

  //Wire declarations for instance 'or_423' (Module coreir_or)
  wire [15:0] or_423__in0;
  wire [15:0] or_423__in1;
  wire [15:0] or_423__out;
  coreir_or #(.width(16)) or_423(
    .in0(or_423__in0),
    .in1(or_423__in1),
    .out(or_423__out)
  );

  //Wire declarations for instance 'or_425' (Module coreir_or)
  wire [15:0] or_425__in0;
  wire [15:0] or_425__in1;
  wire [15:0] or_425__out;
  coreir_or #(.width(16)) or_425(
    .in0(or_425__in0),
    .in1(or_425__in1),
    .out(or_425__out)
  );

  //Wire declarations for instance 'or_427' (Module coreir_or)
  wire [15:0] or_427__in0;
  wire [15:0] or_427__in1;
  wire [15:0] or_427__out;
  coreir_or #(.width(16)) or_427(
    .in0(or_427__in0),
    .in1(or_427__in1),
    .out(or_427__out)
  );

  //Wire declarations for instance 'or_429' (Module coreir_or)
  wire [15:0] or_429__in0;
  wire [15:0] or_429__in1;
  wire [15:0] or_429__out;
  coreir_or #(.width(16)) or_429(
    .in0(or_429__in0),
    .in1(or_429__in1),
    .out(or_429__out)
  );

  //Wire declarations for instance 'or_43' (Module coreir_or)
  wire [15:0] or_43__in0;
  wire [15:0] or_43__in1;
  wire [15:0] or_43__out;
  coreir_or #(.width(16)) or_43(
    .in0(or_43__in0),
    .in1(or_43__in1),
    .out(or_43__out)
  );

  //Wire declarations for instance 'or_431' (Module coreir_or)
  wire [15:0] or_431__in0;
  wire [15:0] or_431__in1;
  wire [15:0] or_431__out;
  coreir_or #(.width(16)) or_431(
    .in0(or_431__in0),
    .in1(or_431__in1),
    .out(or_431__out)
  );

  //Wire declarations for instance 'or_433' (Module coreir_or)
  wire [15:0] or_433__in0;
  wire [15:0] or_433__in1;
  wire [15:0] or_433__out;
  coreir_or #(.width(16)) or_433(
    .in0(or_433__in0),
    .in1(or_433__in1),
    .out(or_433__out)
  );

  //Wire declarations for instance 'or_435' (Module coreir_or)
  wire [15:0] or_435__in0;
  wire [15:0] or_435__in1;
  wire [15:0] or_435__out;
  coreir_or #(.width(16)) or_435(
    .in0(or_435__in0),
    .in1(or_435__in1),
    .out(or_435__out)
  );

  //Wire declarations for instance 'or_437' (Module coreir_or)
  wire [15:0] or_437__in0;
  wire [15:0] or_437__in1;
  wire [15:0] or_437__out;
  coreir_or #(.width(16)) or_437(
    .in0(or_437__in0),
    .in1(or_437__in1),
    .out(or_437__out)
  );

  //Wire declarations for instance 'or_439' (Module coreir_or)
  wire [15:0] or_439__in0;
  wire [15:0] or_439__in1;
  wire [15:0] or_439__out;
  coreir_or #(.width(16)) or_439(
    .in0(or_439__in0),
    .in1(or_439__in1),
    .out(or_439__out)
  );

  //Wire declarations for instance 'or_441' (Module coreir_or)
  wire [15:0] or_441__in0;
  wire [15:0] or_441__in1;
  wire [15:0] or_441__out;
  coreir_or #(.width(16)) or_441(
    .in0(or_441__in0),
    .in1(or_441__in1),
    .out(or_441__out)
  );

  //Wire declarations for instance 'or_443' (Module coreir_or)
  wire [15:0] or_443__in0;
  wire [15:0] or_443__in1;
  wire [15:0] or_443__out;
  coreir_or #(.width(16)) or_443(
    .in0(or_443__in0),
    .in1(or_443__in1),
    .out(or_443__out)
  );

  //Wire declarations for instance 'or_445' (Module coreir_or)
  wire [15:0] or_445__in0;
  wire [15:0] or_445__in1;
  wire [15:0] or_445__out;
  coreir_or #(.width(16)) or_445(
    .in0(or_445__in0),
    .in1(or_445__in1),
    .out(or_445__out)
  );

  //Wire declarations for instance 'or_447' (Module coreir_or)
  wire [15:0] or_447__in0;
  wire [15:0] or_447__in1;
  wire [15:0] or_447__out;
  coreir_or #(.width(16)) or_447(
    .in0(or_447__in0),
    .in1(or_447__in1),
    .out(or_447__out)
  );

  //Wire declarations for instance 'or_449' (Module coreir_or)
  wire [15:0] or_449__in0;
  wire [15:0] or_449__in1;
  wire [15:0] or_449__out;
  coreir_or #(.width(16)) or_449(
    .in0(or_449__in0),
    .in1(or_449__in1),
    .out(or_449__out)
  );

  //Wire declarations for instance 'or_45' (Module coreir_or)
  wire [15:0] or_45__in0;
  wire [15:0] or_45__in1;
  wire [15:0] or_45__out;
  coreir_or #(.width(16)) or_45(
    .in0(or_45__in0),
    .in1(or_45__in1),
    .out(or_45__out)
  );

  //Wire declarations for instance 'or_451' (Module coreir_or)
  wire [15:0] or_451__in0;
  wire [15:0] or_451__in1;
  wire [15:0] or_451__out;
  coreir_or #(.width(16)) or_451(
    .in0(or_451__in0),
    .in1(or_451__in1),
    .out(or_451__out)
  );

  //Wire declarations for instance 'or_453' (Module coreir_or)
  wire [15:0] or_453__in0;
  wire [15:0] or_453__in1;
  wire [15:0] or_453__out;
  coreir_or #(.width(16)) or_453(
    .in0(or_453__in0),
    .in1(or_453__in1),
    .out(or_453__out)
  );

  //Wire declarations for instance 'or_455' (Module coreir_or)
  wire [15:0] or_455__in0;
  wire [15:0] or_455__in1;
  wire [15:0] or_455__out;
  coreir_or #(.width(16)) or_455(
    .in0(or_455__in0),
    .in1(or_455__in1),
    .out(or_455__out)
  );

  //Wire declarations for instance 'or_457' (Module coreir_or)
  wire [15:0] or_457__in0;
  wire [15:0] or_457__in1;
  wire [15:0] or_457__out;
  coreir_or #(.width(16)) or_457(
    .in0(or_457__in0),
    .in1(or_457__in1),
    .out(or_457__out)
  );

  //Wire declarations for instance 'or_459' (Module coreir_or)
  wire [15:0] or_459__in0;
  wire [15:0] or_459__in1;
  wire [15:0] or_459__out;
  coreir_or #(.width(16)) or_459(
    .in0(or_459__in0),
    .in1(or_459__in1),
    .out(or_459__out)
  );

  //Wire declarations for instance 'or_461' (Module coreir_or)
  wire [15:0] or_461__in0;
  wire [15:0] or_461__in1;
  wire [15:0] or_461__out;
  coreir_or #(.width(16)) or_461(
    .in0(or_461__in0),
    .in1(or_461__in1),
    .out(or_461__out)
  );

  //Wire declarations for instance 'or_463' (Module coreir_or)
  wire [15:0] or_463__in0;
  wire [15:0] or_463__in1;
  wire [15:0] or_463__out;
  coreir_or #(.width(16)) or_463(
    .in0(or_463__in0),
    .in1(or_463__in1),
    .out(or_463__out)
  );

  //Wire declarations for instance 'or_465' (Module coreir_or)
  wire [15:0] or_465__in0;
  wire [15:0] or_465__in1;
  wire [15:0] or_465__out;
  coreir_or #(.width(16)) or_465(
    .in0(or_465__in0),
    .in1(or_465__in1),
    .out(or_465__out)
  );

  //Wire declarations for instance 'or_467' (Module coreir_or)
  wire [15:0] or_467__in0;
  wire [15:0] or_467__in1;
  wire [15:0] or_467__out;
  coreir_or #(.width(16)) or_467(
    .in0(or_467__in0),
    .in1(or_467__in1),
    .out(or_467__out)
  );

  //Wire declarations for instance 'or_469' (Module coreir_or)
  wire [15:0] or_469__in0;
  wire [15:0] or_469__in1;
  wire [15:0] or_469__out;
  coreir_or #(.width(16)) or_469(
    .in0(or_469__in0),
    .in1(or_469__in1),
    .out(or_469__out)
  );

  //Wire declarations for instance 'or_47' (Module coreir_or)
  wire [15:0] or_47__in0;
  wire [15:0] or_47__in1;
  wire [15:0] or_47__out;
  coreir_or #(.width(16)) or_47(
    .in0(or_47__in0),
    .in1(or_47__in1),
    .out(or_47__out)
  );

  //Wire declarations for instance 'or_471' (Module coreir_or)
  wire [15:0] or_471__in0;
  wire [15:0] or_471__in1;
  wire [15:0] or_471__out;
  coreir_or #(.width(16)) or_471(
    .in0(or_471__in0),
    .in1(or_471__in1),
    .out(or_471__out)
  );

  //Wire declarations for instance 'or_473' (Module coreir_or)
  wire [15:0] or_473__in0;
  wire [15:0] or_473__in1;
  wire [15:0] or_473__out;
  coreir_or #(.width(16)) or_473(
    .in0(or_473__in0),
    .in1(or_473__in1),
    .out(or_473__out)
  );

  //Wire declarations for instance 'or_475' (Module coreir_or)
  wire [15:0] or_475__in0;
  wire [15:0] or_475__in1;
  wire [15:0] or_475__out;
  coreir_or #(.width(16)) or_475(
    .in0(or_475__in0),
    .in1(or_475__in1),
    .out(or_475__out)
  );

  //Wire declarations for instance 'or_477' (Module coreir_or)
  wire [15:0] or_477__in0;
  wire [15:0] or_477__in1;
  wire [15:0] or_477__out;
  coreir_or #(.width(16)) or_477(
    .in0(or_477__in0),
    .in1(or_477__in1),
    .out(or_477__out)
  );

  //Wire declarations for instance 'or_479' (Module coreir_or)
  wire [15:0] or_479__in0;
  wire [15:0] or_479__in1;
  wire [15:0] or_479__out;
  coreir_or #(.width(16)) or_479(
    .in0(or_479__in0),
    .in1(or_479__in1),
    .out(or_479__out)
  );

  //Wire declarations for instance 'or_481' (Module coreir_or)
  wire [15:0] or_481__in0;
  wire [15:0] or_481__in1;
  wire [15:0] or_481__out;
  coreir_or #(.width(16)) or_481(
    .in0(or_481__in0),
    .in1(or_481__in1),
    .out(or_481__out)
  );

  //Wire declarations for instance 'or_483' (Module coreir_or)
  wire [15:0] or_483__in0;
  wire [15:0] or_483__in1;
  wire [15:0] or_483__out;
  coreir_or #(.width(16)) or_483(
    .in0(or_483__in0),
    .in1(or_483__in1),
    .out(or_483__out)
  );

  //Wire declarations for instance 'or_485' (Module coreir_or)
  wire [15:0] or_485__in0;
  wire [15:0] or_485__in1;
  wire [15:0] or_485__out;
  coreir_or #(.width(16)) or_485(
    .in0(or_485__in0),
    .in1(or_485__in1),
    .out(or_485__out)
  );

  //Wire declarations for instance 'or_487' (Module coreir_or)
  wire [15:0] or_487__in0;
  wire [15:0] or_487__in1;
  wire [15:0] or_487__out;
  coreir_or #(.width(16)) or_487(
    .in0(or_487__in0),
    .in1(or_487__in1),
    .out(or_487__out)
  );

  //Wire declarations for instance 'or_489' (Module coreir_or)
  wire [15:0] or_489__in0;
  wire [15:0] or_489__in1;
  wire [15:0] or_489__out;
  coreir_or #(.width(16)) or_489(
    .in0(or_489__in0),
    .in1(or_489__in1),
    .out(or_489__out)
  );

  //Wire declarations for instance 'or_49' (Module coreir_or)
  wire [15:0] or_49__in0;
  wire [15:0] or_49__in1;
  wire [15:0] or_49__out;
  coreir_or #(.width(16)) or_49(
    .in0(or_49__in0),
    .in1(or_49__in1),
    .out(or_49__out)
  );

  //Wire declarations for instance 'or_491' (Module coreir_or)
  wire [15:0] or_491__in0;
  wire [15:0] or_491__in1;
  wire [15:0] or_491__out;
  coreir_or #(.width(16)) or_491(
    .in0(or_491__in0),
    .in1(or_491__in1),
    .out(or_491__out)
  );

  //Wire declarations for instance 'or_493' (Module coreir_or)
  wire [15:0] or_493__in0;
  wire [15:0] or_493__in1;
  wire [15:0] or_493__out;
  coreir_or #(.width(16)) or_493(
    .in0(or_493__in0),
    .in1(or_493__in1),
    .out(or_493__out)
  );

  //Wire declarations for instance 'or_495' (Module coreir_or)
  wire [15:0] or_495__in0;
  wire [15:0] or_495__in1;
  wire [15:0] or_495__out;
  coreir_or #(.width(16)) or_495(
    .in0(or_495__in0),
    .in1(or_495__in1),
    .out(or_495__out)
  );

  //Wire declarations for instance 'or_497' (Module coreir_or)
  wire [15:0] or_497__in0;
  wire [15:0] or_497__in1;
  wire [15:0] or_497__out;
  coreir_or #(.width(16)) or_497(
    .in0(or_497__in0),
    .in1(or_497__in1),
    .out(or_497__out)
  );

  //Wire declarations for instance 'or_499' (Module coreir_or)
  wire [15:0] or_499__in0;
  wire [15:0] or_499__in1;
  wire [15:0] or_499__out;
  coreir_or #(.width(16)) or_499(
    .in0(or_499__in0),
    .in1(or_499__in1),
    .out(or_499__out)
  );

  //Wire declarations for instance 'or_5' (Module coreir_or)
  wire [15:0] or_5__in0;
  wire [15:0] or_5__in1;
  wire [15:0] or_5__out;
  coreir_or #(.width(16)) or_5(
    .in0(or_5__in0),
    .in1(or_5__in1),
    .out(or_5__out)
  );

  //Wire declarations for instance 'or_501' (Module coreir_or)
  wire [15:0] or_501__in0;
  wire [15:0] or_501__in1;
  wire [15:0] or_501__out;
  coreir_or #(.width(16)) or_501(
    .in0(or_501__in0),
    .in1(or_501__in1),
    .out(or_501__out)
  );

  //Wire declarations for instance 'or_503' (Module coreir_or)
  wire [15:0] or_503__in0;
  wire [15:0] or_503__in1;
  wire [15:0] or_503__out;
  coreir_or #(.width(16)) or_503(
    .in0(or_503__in0),
    .in1(or_503__in1),
    .out(or_503__out)
  );

  //Wire declarations for instance 'or_505' (Module coreir_or)
  wire [15:0] or_505__in0;
  wire [15:0] or_505__in1;
  wire [15:0] or_505__out;
  coreir_or #(.width(16)) or_505(
    .in0(or_505__in0),
    .in1(or_505__in1),
    .out(or_505__out)
  );

  //Wire declarations for instance 'or_507' (Module coreir_or)
  wire [15:0] or_507__in0;
  wire [15:0] or_507__in1;
  wire [15:0] or_507__out;
  coreir_or #(.width(16)) or_507(
    .in0(or_507__in0),
    .in1(or_507__in1),
    .out(or_507__out)
  );

  //Wire declarations for instance 'or_509' (Module coreir_or)
  wire [15:0] or_509__in0;
  wire [15:0] or_509__in1;
  wire [15:0] or_509__out;
  coreir_or #(.width(16)) or_509(
    .in0(or_509__in0),
    .in1(or_509__in1),
    .out(or_509__out)
  );

  //Wire declarations for instance 'or_51' (Module coreir_or)
  wire [15:0] or_51__in0;
  wire [15:0] or_51__in1;
  wire [15:0] or_51__out;
  coreir_or #(.width(16)) or_51(
    .in0(or_51__in0),
    .in1(or_51__in1),
    .out(or_51__out)
  );

  //Wire declarations for instance 'or_511' (Module coreir_or)
  wire [15:0] or_511__in0;
  wire [15:0] or_511__in1;
  wire [15:0] or_511__out;
  coreir_or #(.width(16)) or_511(
    .in0(or_511__in0),
    .in1(or_511__in1),
    .out(or_511__out)
  );

  //Wire declarations for instance 'or_513' (Module coreir_or)
  wire [15:0] or_513__in0;
  wire [15:0] or_513__in1;
  wire [15:0] or_513__out;
  coreir_or #(.width(16)) or_513(
    .in0(or_513__in0),
    .in1(or_513__in1),
    .out(or_513__out)
  );

  //Wire declarations for instance 'or_515' (Module coreir_or)
  wire [15:0] or_515__in0;
  wire [15:0] or_515__in1;
  wire [15:0] or_515__out;
  coreir_or #(.width(16)) or_515(
    .in0(or_515__in0),
    .in1(or_515__in1),
    .out(or_515__out)
  );

  //Wire declarations for instance 'or_517' (Module coreir_or)
  wire [15:0] or_517__in0;
  wire [15:0] or_517__in1;
  wire [15:0] or_517__out;
  coreir_or #(.width(16)) or_517(
    .in0(or_517__in0),
    .in1(or_517__in1),
    .out(or_517__out)
  );

  //Wire declarations for instance 'or_519' (Module coreir_or)
  wire [15:0] or_519__in0;
  wire [15:0] or_519__in1;
  wire [15:0] or_519__out;
  coreir_or #(.width(16)) or_519(
    .in0(or_519__in0),
    .in1(or_519__in1),
    .out(or_519__out)
  );

  //Wire declarations for instance 'or_521' (Module coreir_or)
  wire [15:0] or_521__in0;
  wire [15:0] or_521__in1;
  wire [15:0] or_521__out;
  coreir_or #(.width(16)) or_521(
    .in0(or_521__in0),
    .in1(or_521__in1),
    .out(or_521__out)
  );

  //Wire declarations for instance 'or_523' (Module coreir_or)
  wire [15:0] or_523__in0;
  wire [15:0] or_523__in1;
  wire [15:0] or_523__out;
  coreir_or #(.width(16)) or_523(
    .in0(or_523__in0),
    .in1(or_523__in1),
    .out(or_523__out)
  );

  //Wire declarations for instance 'or_525' (Module coreir_or)
  wire [15:0] or_525__in0;
  wire [15:0] or_525__in1;
  wire [15:0] or_525__out;
  coreir_or #(.width(16)) or_525(
    .in0(or_525__in0),
    .in1(or_525__in1),
    .out(or_525__out)
  );

  //Wire declarations for instance 'or_527' (Module coreir_or)
  wire [15:0] or_527__in0;
  wire [15:0] or_527__in1;
  wire [15:0] or_527__out;
  coreir_or #(.width(16)) or_527(
    .in0(or_527__in0),
    .in1(or_527__in1),
    .out(or_527__out)
  );

  //Wire declarations for instance 'or_529' (Module coreir_or)
  wire [15:0] or_529__in0;
  wire [15:0] or_529__in1;
  wire [15:0] or_529__out;
  coreir_or #(.width(16)) or_529(
    .in0(or_529__in0),
    .in1(or_529__in1),
    .out(or_529__out)
  );

  //Wire declarations for instance 'or_53' (Module coreir_or)
  wire [15:0] or_53__in0;
  wire [15:0] or_53__in1;
  wire [15:0] or_53__out;
  coreir_or #(.width(16)) or_53(
    .in0(or_53__in0),
    .in1(or_53__in1),
    .out(or_53__out)
  );

  //Wire declarations for instance 'or_531' (Module coreir_or)
  wire [15:0] or_531__in0;
  wire [15:0] or_531__in1;
  wire [15:0] or_531__out;
  coreir_or #(.width(16)) or_531(
    .in0(or_531__in0),
    .in1(or_531__in1),
    .out(or_531__out)
  );

  //Wire declarations for instance 'or_533' (Module coreir_or)
  wire [15:0] or_533__in0;
  wire [15:0] or_533__in1;
  wire [15:0] or_533__out;
  coreir_or #(.width(16)) or_533(
    .in0(or_533__in0),
    .in1(or_533__in1),
    .out(or_533__out)
  );

  //Wire declarations for instance 'or_535' (Module coreir_or)
  wire [15:0] or_535__in0;
  wire [15:0] or_535__in1;
  wire [15:0] or_535__out;
  coreir_or #(.width(16)) or_535(
    .in0(or_535__in0),
    .in1(or_535__in1),
    .out(or_535__out)
  );

  //Wire declarations for instance 'or_537' (Module coreir_or)
  wire [15:0] or_537__in0;
  wire [15:0] or_537__in1;
  wire [15:0] or_537__out;
  coreir_or #(.width(16)) or_537(
    .in0(or_537__in0),
    .in1(or_537__in1),
    .out(or_537__out)
  );

  //Wire declarations for instance 'or_539' (Module coreir_or)
  wire [15:0] or_539__in0;
  wire [15:0] or_539__in1;
  wire [15:0] or_539__out;
  coreir_or #(.width(16)) or_539(
    .in0(or_539__in0),
    .in1(or_539__in1),
    .out(or_539__out)
  );

  //Wire declarations for instance 'or_541' (Module coreir_or)
  wire [15:0] or_541__in0;
  wire [15:0] or_541__in1;
  wire [15:0] or_541__out;
  coreir_or #(.width(16)) or_541(
    .in0(or_541__in0),
    .in1(or_541__in1),
    .out(or_541__out)
  );

  //Wire declarations for instance 'or_543' (Module coreir_or)
  wire [15:0] or_543__in0;
  wire [15:0] or_543__in1;
  wire [15:0] or_543__out;
  coreir_or #(.width(16)) or_543(
    .in0(or_543__in0),
    .in1(or_543__in1),
    .out(or_543__out)
  );

  //Wire declarations for instance 'or_545' (Module coreir_or)
  wire [15:0] or_545__in0;
  wire [15:0] or_545__in1;
  wire [15:0] or_545__out;
  coreir_or #(.width(16)) or_545(
    .in0(or_545__in0),
    .in1(or_545__in1),
    .out(or_545__out)
  );

  //Wire declarations for instance 'or_547' (Module coreir_or)
  wire [15:0] or_547__in0;
  wire [15:0] or_547__in1;
  wire [15:0] or_547__out;
  coreir_or #(.width(16)) or_547(
    .in0(or_547__in0),
    .in1(or_547__in1),
    .out(or_547__out)
  );

  //Wire declarations for instance 'or_549' (Module coreir_or)
  wire [15:0] or_549__in0;
  wire [15:0] or_549__in1;
  wire [15:0] or_549__out;
  coreir_or #(.width(16)) or_549(
    .in0(or_549__in0),
    .in1(or_549__in1),
    .out(or_549__out)
  );

  //Wire declarations for instance 'or_55' (Module coreir_or)
  wire [15:0] or_55__in0;
  wire [15:0] or_55__in1;
  wire [15:0] or_55__out;
  coreir_or #(.width(16)) or_55(
    .in0(or_55__in0),
    .in1(or_55__in1),
    .out(or_55__out)
  );

  //Wire declarations for instance 'or_551' (Module coreir_or)
  wire [15:0] or_551__in0;
  wire [15:0] or_551__in1;
  wire [15:0] or_551__out;
  coreir_or #(.width(16)) or_551(
    .in0(or_551__in0),
    .in1(or_551__in1),
    .out(or_551__out)
  );

  //Wire declarations for instance 'or_553' (Module coreir_or)
  wire [15:0] or_553__in0;
  wire [15:0] or_553__in1;
  wire [15:0] or_553__out;
  coreir_or #(.width(16)) or_553(
    .in0(or_553__in0),
    .in1(or_553__in1),
    .out(or_553__out)
  );

  //Wire declarations for instance 'or_555' (Module coreir_or)
  wire [15:0] or_555__in0;
  wire [15:0] or_555__in1;
  wire [15:0] or_555__out;
  coreir_or #(.width(16)) or_555(
    .in0(or_555__in0),
    .in1(or_555__in1),
    .out(or_555__out)
  );

  //Wire declarations for instance 'or_557' (Module coreir_or)
  wire [15:0] or_557__in0;
  wire [15:0] or_557__in1;
  wire [15:0] or_557__out;
  coreir_or #(.width(16)) or_557(
    .in0(or_557__in0),
    .in1(or_557__in1),
    .out(or_557__out)
  );

  //Wire declarations for instance 'or_559' (Module coreir_or)
  wire [15:0] or_559__in0;
  wire [15:0] or_559__in1;
  wire [15:0] or_559__out;
  coreir_or #(.width(16)) or_559(
    .in0(or_559__in0),
    .in1(or_559__in1),
    .out(or_559__out)
  );

  //Wire declarations for instance 'or_561' (Module coreir_or)
  wire [15:0] or_561__in0;
  wire [15:0] or_561__in1;
  wire [15:0] or_561__out;
  coreir_or #(.width(16)) or_561(
    .in0(or_561__in0),
    .in1(or_561__in1),
    .out(or_561__out)
  );

  //Wire declarations for instance 'or_563' (Module coreir_or)
  wire [15:0] or_563__in0;
  wire [15:0] or_563__in1;
  wire [15:0] or_563__out;
  coreir_or #(.width(16)) or_563(
    .in0(or_563__in0),
    .in1(or_563__in1),
    .out(or_563__out)
  );

  //Wire declarations for instance 'or_565' (Module coreir_or)
  wire [15:0] or_565__in0;
  wire [15:0] or_565__in1;
  wire [15:0] or_565__out;
  coreir_or #(.width(16)) or_565(
    .in0(or_565__in0),
    .in1(or_565__in1),
    .out(or_565__out)
  );

  //Wire declarations for instance 'or_567' (Module coreir_or)
  wire [15:0] or_567__in0;
  wire [15:0] or_567__in1;
  wire [15:0] or_567__out;
  coreir_or #(.width(16)) or_567(
    .in0(or_567__in0),
    .in1(or_567__in1),
    .out(or_567__out)
  );

  //Wire declarations for instance 'or_569' (Module coreir_or)
  wire [15:0] or_569__in0;
  wire [15:0] or_569__in1;
  wire [15:0] or_569__out;
  coreir_or #(.width(16)) or_569(
    .in0(or_569__in0),
    .in1(or_569__in1),
    .out(or_569__out)
  );

  //Wire declarations for instance 'or_57' (Module coreir_or)
  wire [15:0] or_57__in0;
  wire [15:0] or_57__in1;
  wire [15:0] or_57__out;
  coreir_or #(.width(16)) or_57(
    .in0(or_57__in0),
    .in1(or_57__in1),
    .out(or_57__out)
  );

  //Wire declarations for instance 'or_571' (Module coreir_or)
  wire [15:0] or_571__in0;
  wire [15:0] or_571__in1;
  wire [15:0] or_571__out;
  coreir_or #(.width(16)) or_571(
    .in0(or_571__in0),
    .in1(or_571__in1),
    .out(or_571__out)
  );

  //Wire declarations for instance 'or_573' (Module coreir_or)
  wire [15:0] or_573__in0;
  wire [15:0] or_573__in1;
  wire [15:0] or_573__out;
  coreir_or #(.width(16)) or_573(
    .in0(or_573__in0),
    .in1(or_573__in1),
    .out(or_573__out)
  );

  //Wire declarations for instance 'or_575' (Module coreir_or)
  wire [15:0] or_575__in0;
  wire [15:0] or_575__in1;
  wire [15:0] or_575__out;
  coreir_or #(.width(16)) or_575(
    .in0(or_575__in0),
    .in1(or_575__in1),
    .out(or_575__out)
  );

  //Wire declarations for instance 'or_577' (Module coreir_or)
  wire [15:0] or_577__in0;
  wire [15:0] or_577__in1;
  wire [15:0] or_577__out;
  coreir_or #(.width(16)) or_577(
    .in0(or_577__in0),
    .in1(or_577__in1),
    .out(or_577__out)
  );

  //Wire declarations for instance 'or_579' (Module coreir_or)
  wire [15:0] or_579__in0;
  wire [15:0] or_579__in1;
  wire [15:0] or_579__out;
  coreir_or #(.width(16)) or_579(
    .in0(or_579__in0),
    .in1(or_579__in1),
    .out(or_579__out)
  );

  //Wire declarations for instance 'or_581' (Module coreir_or)
  wire [15:0] or_581__in0;
  wire [15:0] or_581__in1;
  wire [15:0] or_581__out;
  coreir_or #(.width(16)) or_581(
    .in0(or_581__in0),
    .in1(or_581__in1),
    .out(or_581__out)
  );

  //Wire declarations for instance 'or_583' (Module coreir_or)
  wire [15:0] or_583__in0;
  wire [15:0] or_583__in1;
  wire [15:0] or_583__out;
  coreir_or #(.width(16)) or_583(
    .in0(or_583__in0),
    .in1(or_583__in1),
    .out(or_583__out)
  );

  //Wire declarations for instance 'or_585' (Module coreir_or)
  wire [15:0] or_585__in0;
  wire [15:0] or_585__in1;
  wire [15:0] or_585__out;
  coreir_or #(.width(16)) or_585(
    .in0(or_585__in0),
    .in1(or_585__in1),
    .out(or_585__out)
  );

  //Wire declarations for instance 'or_587' (Module coreir_or)
  wire [15:0] or_587__in0;
  wire [15:0] or_587__in1;
  wire [15:0] or_587__out;
  coreir_or #(.width(16)) or_587(
    .in0(or_587__in0),
    .in1(or_587__in1),
    .out(or_587__out)
  );

  //Wire declarations for instance 'or_589' (Module coreir_or)
  wire [15:0] or_589__in0;
  wire [15:0] or_589__in1;
  wire [15:0] or_589__out;
  coreir_or #(.width(16)) or_589(
    .in0(or_589__in0),
    .in1(or_589__in1),
    .out(or_589__out)
  );

  //Wire declarations for instance 'or_59' (Module coreir_or)
  wire [15:0] or_59__in0;
  wire [15:0] or_59__in1;
  wire [15:0] or_59__out;
  coreir_or #(.width(16)) or_59(
    .in0(or_59__in0),
    .in1(or_59__in1),
    .out(or_59__out)
  );

  //Wire declarations for instance 'or_591' (Module coreir_or)
  wire [15:0] or_591__in0;
  wire [15:0] or_591__in1;
  wire [15:0] or_591__out;
  coreir_or #(.width(16)) or_591(
    .in0(or_591__in0),
    .in1(or_591__in1),
    .out(or_591__out)
  );

  //Wire declarations for instance 'or_593' (Module coreir_or)
  wire [15:0] or_593__in0;
  wire [15:0] or_593__in1;
  wire [15:0] or_593__out;
  coreir_or #(.width(16)) or_593(
    .in0(or_593__in0),
    .in1(or_593__in1),
    .out(or_593__out)
  );

  //Wire declarations for instance 'or_595' (Module coreir_or)
  wire [15:0] or_595__in0;
  wire [15:0] or_595__in1;
  wire [15:0] or_595__out;
  coreir_or #(.width(16)) or_595(
    .in0(or_595__in0),
    .in1(or_595__in1),
    .out(or_595__out)
  );

  //Wire declarations for instance 'or_597' (Module coreir_or)
  wire [15:0] or_597__in0;
  wire [15:0] or_597__in1;
  wire [15:0] or_597__out;
  coreir_or #(.width(16)) or_597(
    .in0(or_597__in0),
    .in1(or_597__in1),
    .out(or_597__out)
  );

  //Wire declarations for instance 'or_599' (Module coreir_or)
  wire [15:0] or_599__in0;
  wire [15:0] or_599__in1;
  wire [15:0] or_599__out;
  coreir_or #(.width(16)) or_599(
    .in0(or_599__in0),
    .in1(or_599__in1),
    .out(or_599__out)
  );

  //Wire declarations for instance 'or_601' (Module coreir_or)
  wire [15:0] or_601__in0;
  wire [15:0] or_601__in1;
  wire [15:0] or_601__out;
  coreir_or #(.width(16)) or_601(
    .in0(or_601__in0),
    .in1(or_601__in1),
    .out(or_601__out)
  );

  //Wire declarations for instance 'or_603' (Module coreir_or)
  wire [15:0] or_603__in0;
  wire [15:0] or_603__in1;
  wire [15:0] or_603__out;
  coreir_or #(.width(16)) or_603(
    .in0(or_603__in0),
    .in1(or_603__in1),
    .out(or_603__out)
  );

  //Wire declarations for instance 'or_605' (Module coreir_or)
  wire [15:0] or_605__in0;
  wire [15:0] or_605__in1;
  wire [15:0] or_605__out;
  coreir_or #(.width(16)) or_605(
    .in0(or_605__in0),
    .in1(or_605__in1),
    .out(or_605__out)
  );

  //Wire declarations for instance 'or_607' (Module coreir_or)
  wire [15:0] or_607__in0;
  wire [15:0] or_607__in1;
  wire [15:0] or_607__out;
  coreir_or #(.width(16)) or_607(
    .in0(or_607__in0),
    .in1(or_607__in1),
    .out(or_607__out)
  );

  //Wire declarations for instance 'or_609' (Module coreir_or)
  wire [15:0] or_609__in0;
  wire [15:0] or_609__in1;
  wire [15:0] or_609__out;
  coreir_or #(.width(16)) or_609(
    .in0(or_609__in0),
    .in1(or_609__in1),
    .out(or_609__out)
  );

  //Wire declarations for instance 'or_61' (Module coreir_or)
  wire [15:0] or_61__in0;
  wire [15:0] or_61__in1;
  wire [15:0] or_61__out;
  coreir_or #(.width(16)) or_61(
    .in0(or_61__in0),
    .in1(or_61__in1),
    .out(or_61__out)
  );

  //Wire declarations for instance 'or_611' (Module coreir_or)
  wire [15:0] or_611__in0;
  wire [15:0] or_611__in1;
  wire [15:0] or_611__out;
  coreir_or #(.width(16)) or_611(
    .in0(or_611__in0),
    .in1(or_611__in1),
    .out(or_611__out)
  );

  //Wire declarations for instance 'or_613' (Module coreir_or)
  wire [15:0] or_613__in0;
  wire [15:0] or_613__in1;
  wire [15:0] or_613__out;
  coreir_or #(.width(16)) or_613(
    .in0(or_613__in0),
    .in1(or_613__in1),
    .out(or_613__out)
  );

  //Wire declarations for instance 'or_615' (Module coreir_or)
  wire [15:0] or_615__in0;
  wire [15:0] or_615__in1;
  wire [15:0] or_615__out;
  coreir_or #(.width(16)) or_615(
    .in0(or_615__in0),
    .in1(or_615__in1),
    .out(or_615__out)
  );

  //Wire declarations for instance 'or_617' (Module coreir_or)
  wire [15:0] or_617__in0;
  wire [15:0] or_617__in1;
  wire [15:0] or_617__out;
  coreir_or #(.width(16)) or_617(
    .in0(or_617__in0),
    .in1(or_617__in1),
    .out(or_617__out)
  );

  //Wire declarations for instance 'or_619' (Module coreir_or)
  wire [15:0] or_619__in0;
  wire [15:0] or_619__in1;
  wire [15:0] or_619__out;
  coreir_or #(.width(16)) or_619(
    .in0(or_619__in0),
    .in1(or_619__in1),
    .out(or_619__out)
  );

  //Wire declarations for instance 'or_621' (Module coreir_or)
  wire [15:0] or_621__in0;
  wire [15:0] or_621__in1;
  wire [15:0] or_621__out;
  coreir_or #(.width(16)) or_621(
    .in0(or_621__in0),
    .in1(or_621__in1),
    .out(or_621__out)
  );

  //Wire declarations for instance 'or_623' (Module coreir_or)
  wire [15:0] or_623__in0;
  wire [15:0] or_623__in1;
  wire [15:0] or_623__out;
  coreir_or #(.width(16)) or_623(
    .in0(or_623__in0),
    .in1(or_623__in1),
    .out(or_623__out)
  );

  //Wire declarations for instance 'or_625' (Module coreir_or)
  wire [15:0] or_625__in0;
  wire [15:0] or_625__in1;
  wire [15:0] or_625__out;
  coreir_or #(.width(16)) or_625(
    .in0(or_625__in0),
    .in1(or_625__in1),
    .out(or_625__out)
  );

  //Wire declarations for instance 'or_627' (Module coreir_or)
  wire [15:0] or_627__in0;
  wire [15:0] or_627__in1;
  wire [15:0] or_627__out;
  coreir_or #(.width(16)) or_627(
    .in0(or_627__in0),
    .in1(or_627__in1),
    .out(or_627__out)
  );

  //Wire declarations for instance 'or_629' (Module coreir_or)
  wire [15:0] or_629__in0;
  wire [15:0] or_629__in1;
  wire [15:0] or_629__out;
  coreir_or #(.width(16)) or_629(
    .in0(or_629__in0),
    .in1(or_629__in1),
    .out(or_629__out)
  );

  //Wire declarations for instance 'or_63' (Module coreir_or)
  wire [15:0] or_63__in0;
  wire [15:0] or_63__in1;
  wire [15:0] or_63__out;
  coreir_or #(.width(16)) or_63(
    .in0(or_63__in0),
    .in1(or_63__in1),
    .out(or_63__out)
  );

  //Wire declarations for instance 'or_631' (Module coreir_or)
  wire [15:0] or_631__in0;
  wire [15:0] or_631__in1;
  wire [15:0] or_631__out;
  coreir_or #(.width(16)) or_631(
    .in0(or_631__in0),
    .in1(or_631__in1),
    .out(or_631__out)
  );

  //Wire declarations for instance 'or_633' (Module coreir_or)
  wire [15:0] or_633__in0;
  wire [15:0] or_633__in1;
  wire [15:0] or_633__out;
  coreir_or #(.width(16)) or_633(
    .in0(or_633__in0),
    .in1(or_633__in1),
    .out(or_633__out)
  );

  //Wire declarations for instance 'or_635' (Module coreir_or)
  wire [15:0] or_635__in0;
  wire [15:0] or_635__in1;
  wire [15:0] or_635__out;
  coreir_or #(.width(16)) or_635(
    .in0(or_635__in0),
    .in1(or_635__in1),
    .out(or_635__out)
  );

  //Wire declarations for instance 'or_637' (Module coreir_or)
  wire [15:0] or_637__in0;
  wire [15:0] or_637__in1;
  wire [15:0] or_637__out;
  coreir_or #(.width(16)) or_637(
    .in0(or_637__in0),
    .in1(or_637__in1),
    .out(or_637__out)
  );

  //Wire declarations for instance 'or_639' (Module coreir_or)
  wire [15:0] or_639__in0;
  wire [15:0] or_639__in1;
  wire [15:0] or_639__out;
  coreir_or #(.width(16)) or_639(
    .in0(or_639__in0),
    .in1(or_639__in1),
    .out(or_639__out)
  );

  //Wire declarations for instance 'or_641' (Module coreir_or)
  wire [15:0] or_641__in0;
  wire [15:0] or_641__in1;
  wire [15:0] or_641__out;
  coreir_or #(.width(16)) or_641(
    .in0(or_641__in0),
    .in1(or_641__in1),
    .out(or_641__out)
  );

  //Wire declarations for instance 'or_643' (Module coreir_or)
  wire [15:0] or_643__in0;
  wire [15:0] or_643__in1;
  wire [15:0] or_643__out;
  coreir_or #(.width(16)) or_643(
    .in0(or_643__in0),
    .in1(or_643__in1),
    .out(or_643__out)
  );

  //Wire declarations for instance 'or_645' (Module coreir_or)
  wire [15:0] or_645__in0;
  wire [15:0] or_645__in1;
  wire [15:0] or_645__out;
  coreir_or #(.width(16)) or_645(
    .in0(or_645__in0),
    .in1(or_645__in1),
    .out(or_645__out)
  );

  //Wire declarations for instance 'or_647' (Module coreir_or)
  wire [15:0] or_647__in0;
  wire [15:0] or_647__in1;
  wire [15:0] or_647__out;
  coreir_or #(.width(16)) or_647(
    .in0(or_647__in0),
    .in1(or_647__in1),
    .out(or_647__out)
  );

  //Wire declarations for instance 'or_649' (Module coreir_or)
  wire [15:0] or_649__in0;
  wire [15:0] or_649__in1;
  wire [15:0] or_649__out;
  coreir_or #(.width(16)) or_649(
    .in0(or_649__in0),
    .in1(or_649__in1),
    .out(or_649__out)
  );

  //Wire declarations for instance 'or_65' (Module coreir_or)
  wire [15:0] or_65__in0;
  wire [15:0] or_65__in1;
  wire [15:0] or_65__out;
  coreir_or #(.width(16)) or_65(
    .in0(or_65__in0),
    .in1(or_65__in1),
    .out(or_65__out)
  );

  //Wire declarations for instance 'or_651' (Module coreir_or)
  wire [15:0] or_651__in0;
  wire [15:0] or_651__in1;
  wire [15:0] or_651__out;
  coreir_or #(.width(16)) or_651(
    .in0(or_651__in0),
    .in1(or_651__in1),
    .out(or_651__out)
  );

  //Wire declarations for instance 'or_653' (Module coreir_or)
  wire [15:0] or_653__in0;
  wire [15:0] or_653__in1;
  wire [15:0] or_653__out;
  coreir_or #(.width(16)) or_653(
    .in0(or_653__in0),
    .in1(or_653__in1),
    .out(or_653__out)
  );

  //Wire declarations for instance 'or_655' (Module coreir_or)
  wire [15:0] or_655__in0;
  wire [15:0] or_655__in1;
  wire [15:0] or_655__out;
  coreir_or #(.width(16)) or_655(
    .in0(or_655__in0),
    .in1(or_655__in1),
    .out(or_655__out)
  );

  //Wire declarations for instance 'or_657' (Module coreir_or)
  wire [15:0] or_657__in0;
  wire [15:0] or_657__in1;
  wire [15:0] or_657__out;
  coreir_or #(.width(16)) or_657(
    .in0(or_657__in0),
    .in1(or_657__in1),
    .out(or_657__out)
  );

  //Wire declarations for instance 'or_659' (Module coreir_or)
  wire [15:0] or_659__in0;
  wire [15:0] or_659__in1;
  wire [15:0] or_659__out;
  coreir_or #(.width(16)) or_659(
    .in0(or_659__in0),
    .in1(or_659__in1),
    .out(or_659__out)
  );

  //Wire declarations for instance 'or_661' (Module coreir_or)
  wire [15:0] or_661__in0;
  wire [15:0] or_661__in1;
  wire [15:0] or_661__out;
  coreir_or #(.width(16)) or_661(
    .in0(or_661__in0),
    .in1(or_661__in1),
    .out(or_661__out)
  );

  //Wire declarations for instance 'or_663' (Module coreir_or)
  wire [15:0] or_663__in0;
  wire [15:0] or_663__in1;
  wire [15:0] or_663__out;
  coreir_or #(.width(16)) or_663(
    .in0(or_663__in0),
    .in1(or_663__in1),
    .out(or_663__out)
  );

  //Wire declarations for instance 'or_665' (Module coreir_or)
  wire [15:0] or_665__in0;
  wire [15:0] or_665__in1;
  wire [15:0] or_665__out;
  coreir_or #(.width(16)) or_665(
    .in0(or_665__in0),
    .in1(or_665__in1),
    .out(or_665__out)
  );

  //Wire declarations for instance 'or_667' (Module coreir_or)
  wire [15:0] or_667__in0;
  wire [15:0] or_667__in1;
  wire [15:0] or_667__out;
  coreir_or #(.width(16)) or_667(
    .in0(or_667__in0),
    .in1(or_667__in1),
    .out(or_667__out)
  );

  //Wire declarations for instance 'or_669' (Module coreir_or)
  wire [15:0] or_669__in0;
  wire [15:0] or_669__in1;
  wire [15:0] or_669__out;
  coreir_or #(.width(16)) or_669(
    .in0(or_669__in0),
    .in1(or_669__in1),
    .out(or_669__out)
  );

  //Wire declarations for instance 'or_67' (Module coreir_or)
  wire [15:0] or_67__in0;
  wire [15:0] or_67__in1;
  wire [15:0] or_67__out;
  coreir_or #(.width(16)) or_67(
    .in0(or_67__in0),
    .in1(or_67__in1),
    .out(or_67__out)
  );

  //Wire declarations for instance 'or_671' (Module coreir_or)
  wire [15:0] or_671__in0;
  wire [15:0] or_671__in1;
  wire [15:0] or_671__out;
  coreir_or #(.width(16)) or_671(
    .in0(or_671__in0),
    .in1(or_671__in1),
    .out(or_671__out)
  );

  //Wire declarations for instance 'or_673' (Module coreir_or)
  wire [15:0] or_673__in0;
  wire [15:0] or_673__in1;
  wire [15:0] or_673__out;
  coreir_or #(.width(16)) or_673(
    .in0(or_673__in0),
    .in1(or_673__in1),
    .out(or_673__out)
  );

  //Wire declarations for instance 'or_675' (Module coreir_or)
  wire [15:0] or_675__in0;
  wire [15:0] or_675__in1;
  wire [15:0] or_675__out;
  coreir_or #(.width(16)) or_675(
    .in0(or_675__in0),
    .in1(or_675__in1),
    .out(or_675__out)
  );

  //Wire declarations for instance 'or_677' (Module coreir_or)
  wire [15:0] or_677__in0;
  wire [15:0] or_677__in1;
  wire [15:0] or_677__out;
  coreir_or #(.width(16)) or_677(
    .in0(or_677__in0),
    .in1(or_677__in1),
    .out(or_677__out)
  );

  //Wire declarations for instance 'or_679' (Module coreir_or)
  wire [15:0] or_679__in0;
  wire [15:0] or_679__in1;
  wire [15:0] or_679__out;
  coreir_or #(.width(16)) or_679(
    .in0(or_679__in0),
    .in1(or_679__in1),
    .out(or_679__out)
  );

  //Wire declarations for instance 'or_681' (Module coreir_or)
  wire [15:0] or_681__in0;
  wire [15:0] or_681__in1;
  wire [15:0] or_681__out;
  coreir_or #(.width(16)) or_681(
    .in0(or_681__in0),
    .in1(or_681__in1),
    .out(or_681__out)
  );

  //Wire declarations for instance 'or_683' (Module coreir_or)
  wire [15:0] or_683__in0;
  wire [15:0] or_683__in1;
  wire [15:0] or_683__out;
  coreir_or #(.width(16)) or_683(
    .in0(or_683__in0),
    .in1(or_683__in1),
    .out(or_683__out)
  );

  //Wire declarations for instance 'or_685' (Module coreir_or)
  wire [15:0] or_685__in0;
  wire [15:0] or_685__in1;
  wire [15:0] or_685__out;
  coreir_or #(.width(16)) or_685(
    .in0(or_685__in0),
    .in1(or_685__in1),
    .out(or_685__out)
  );

  //Wire declarations for instance 'or_687' (Module coreir_or)
  wire [15:0] or_687__in0;
  wire [15:0] or_687__in1;
  wire [15:0] or_687__out;
  coreir_or #(.width(16)) or_687(
    .in0(or_687__in0),
    .in1(or_687__in1),
    .out(or_687__out)
  );

  //Wire declarations for instance 'or_689' (Module coreir_or)
  wire [15:0] or_689__in0;
  wire [15:0] or_689__in1;
  wire [15:0] or_689__out;
  coreir_or #(.width(16)) or_689(
    .in0(or_689__in0),
    .in1(or_689__in1),
    .out(or_689__out)
  );

  //Wire declarations for instance 'or_69' (Module coreir_or)
  wire [15:0] or_69__in0;
  wire [15:0] or_69__in1;
  wire [15:0] or_69__out;
  coreir_or #(.width(16)) or_69(
    .in0(or_69__in0),
    .in1(or_69__in1),
    .out(or_69__out)
  );

  //Wire declarations for instance 'or_691' (Module coreir_or)
  wire [15:0] or_691__in0;
  wire [15:0] or_691__in1;
  wire [15:0] or_691__out;
  coreir_or #(.width(16)) or_691(
    .in0(or_691__in0),
    .in1(or_691__in1),
    .out(or_691__out)
  );

  //Wire declarations for instance 'or_693' (Module coreir_or)
  wire [15:0] or_693__in0;
  wire [15:0] or_693__in1;
  wire [15:0] or_693__out;
  coreir_or #(.width(16)) or_693(
    .in0(or_693__in0),
    .in1(or_693__in1),
    .out(or_693__out)
  );

  //Wire declarations for instance 'or_695' (Module coreir_or)
  wire [15:0] or_695__in0;
  wire [15:0] or_695__in1;
  wire [15:0] or_695__out;
  coreir_or #(.width(16)) or_695(
    .in0(or_695__in0),
    .in1(or_695__in1),
    .out(or_695__out)
  );

  //Wire declarations for instance 'or_697' (Module coreir_or)
  wire [15:0] or_697__in0;
  wire [15:0] or_697__in1;
  wire [15:0] or_697__out;
  coreir_or #(.width(16)) or_697(
    .in0(or_697__in0),
    .in1(or_697__in1),
    .out(or_697__out)
  );

  //Wire declarations for instance 'or_699' (Module coreir_or)
  wire [15:0] or_699__in0;
  wire [15:0] or_699__in1;
  wire [15:0] or_699__out;
  coreir_or #(.width(16)) or_699(
    .in0(or_699__in0),
    .in1(or_699__in1),
    .out(or_699__out)
  );

  //Wire declarations for instance 'or_7' (Module coreir_or)
  wire [15:0] or_7__in0;
  wire [15:0] or_7__in1;
  wire [15:0] or_7__out;
  coreir_or #(.width(16)) or_7(
    .in0(or_7__in0),
    .in1(or_7__in1),
    .out(or_7__out)
  );

  //Wire declarations for instance 'or_701' (Module coreir_or)
  wire [15:0] or_701__in0;
  wire [15:0] or_701__in1;
  wire [15:0] or_701__out;
  coreir_or #(.width(16)) or_701(
    .in0(or_701__in0),
    .in1(or_701__in1),
    .out(or_701__out)
  );

  //Wire declarations for instance 'or_703' (Module coreir_or)
  wire [15:0] or_703__in0;
  wire [15:0] or_703__in1;
  wire [15:0] or_703__out;
  coreir_or #(.width(16)) or_703(
    .in0(or_703__in0),
    .in1(or_703__in1),
    .out(or_703__out)
  );

  //Wire declarations for instance 'or_705' (Module coreir_or)
  wire [15:0] or_705__in0;
  wire [15:0] or_705__in1;
  wire [15:0] or_705__out;
  coreir_or #(.width(16)) or_705(
    .in0(or_705__in0),
    .in1(or_705__in1),
    .out(or_705__out)
  );

  //Wire declarations for instance 'or_707' (Module coreir_or)
  wire [15:0] or_707__in0;
  wire [15:0] or_707__in1;
  wire [15:0] or_707__out;
  coreir_or #(.width(16)) or_707(
    .in0(or_707__in0),
    .in1(or_707__in1),
    .out(or_707__out)
  );

  //Wire declarations for instance 'or_709' (Module coreir_or)
  wire [15:0] or_709__in0;
  wire [15:0] or_709__in1;
  wire [15:0] or_709__out;
  coreir_or #(.width(16)) or_709(
    .in0(or_709__in0),
    .in1(or_709__in1),
    .out(or_709__out)
  );

  //Wire declarations for instance 'or_71' (Module coreir_or)
  wire [15:0] or_71__in0;
  wire [15:0] or_71__in1;
  wire [15:0] or_71__out;
  coreir_or #(.width(16)) or_71(
    .in0(or_71__in0),
    .in1(or_71__in1),
    .out(or_71__out)
  );

  //Wire declarations for instance 'or_711' (Module coreir_or)
  wire [15:0] or_711__in0;
  wire [15:0] or_711__in1;
  wire [15:0] or_711__out;
  coreir_or #(.width(16)) or_711(
    .in0(or_711__in0),
    .in1(or_711__in1),
    .out(or_711__out)
  );

  //Wire declarations for instance 'or_713' (Module coreir_or)
  wire [15:0] or_713__in0;
  wire [15:0] or_713__in1;
  wire [15:0] or_713__out;
  coreir_or #(.width(16)) or_713(
    .in0(or_713__in0),
    .in1(or_713__in1),
    .out(or_713__out)
  );

  //Wire declarations for instance 'or_715' (Module coreir_or)
  wire [15:0] or_715__in0;
  wire [15:0] or_715__in1;
  wire [15:0] or_715__out;
  coreir_or #(.width(16)) or_715(
    .in0(or_715__in0),
    .in1(or_715__in1),
    .out(or_715__out)
  );

  //Wire declarations for instance 'or_717' (Module coreir_or)
  wire [15:0] or_717__in0;
  wire [15:0] or_717__in1;
  wire [15:0] or_717__out;
  coreir_or #(.width(16)) or_717(
    .in0(or_717__in0),
    .in1(or_717__in1),
    .out(or_717__out)
  );

  //Wire declarations for instance 'or_719' (Module coreir_or)
  wire [15:0] or_719__in0;
  wire [15:0] or_719__in1;
  wire [15:0] or_719__out;
  coreir_or #(.width(16)) or_719(
    .in0(or_719__in0),
    .in1(or_719__in1),
    .out(or_719__out)
  );

  //Wire declarations for instance 'or_721' (Module coreir_or)
  wire [15:0] or_721__in0;
  wire [15:0] or_721__in1;
  wire [15:0] or_721__out;
  coreir_or #(.width(16)) or_721(
    .in0(or_721__in0),
    .in1(or_721__in1),
    .out(or_721__out)
  );

  //Wire declarations for instance 'or_723' (Module coreir_or)
  wire [15:0] or_723__in0;
  wire [15:0] or_723__in1;
  wire [15:0] or_723__out;
  coreir_or #(.width(16)) or_723(
    .in0(or_723__in0),
    .in1(or_723__in1),
    .out(or_723__out)
  );

  //Wire declarations for instance 'or_725' (Module coreir_or)
  wire [15:0] or_725__in0;
  wire [15:0] or_725__in1;
  wire [15:0] or_725__out;
  coreir_or #(.width(16)) or_725(
    .in0(or_725__in0),
    .in1(or_725__in1),
    .out(or_725__out)
  );

  //Wire declarations for instance 'or_727' (Module coreir_or)
  wire [15:0] or_727__in0;
  wire [15:0] or_727__in1;
  wire [15:0] or_727__out;
  coreir_or #(.width(16)) or_727(
    .in0(or_727__in0),
    .in1(or_727__in1),
    .out(or_727__out)
  );

  //Wire declarations for instance 'or_729' (Module coreir_or)
  wire [15:0] or_729__in0;
  wire [15:0] or_729__in1;
  wire [15:0] or_729__out;
  coreir_or #(.width(16)) or_729(
    .in0(or_729__in0),
    .in1(or_729__in1),
    .out(or_729__out)
  );

  //Wire declarations for instance 'or_73' (Module coreir_or)
  wire [15:0] or_73__in0;
  wire [15:0] or_73__in1;
  wire [15:0] or_73__out;
  coreir_or #(.width(16)) or_73(
    .in0(or_73__in0),
    .in1(or_73__in1),
    .out(or_73__out)
  );

  //Wire declarations for instance 'or_731' (Module coreir_or)
  wire [15:0] or_731__in0;
  wire [15:0] or_731__in1;
  wire [15:0] or_731__out;
  coreir_or #(.width(16)) or_731(
    .in0(or_731__in0),
    .in1(or_731__in1),
    .out(or_731__out)
  );

  //Wire declarations for instance 'or_733' (Module coreir_or)
  wire [15:0] or_733__in0;
  wire [15:0] or_733__in1;
  wire [15:0] or_733__out;
  coreir_or #(.width(16)) or_733(
    .in0(or_733__in0),
    .in1(or_733__in1),
    .out(or_733__out)
  );

  //Wire declarations for instance 'or_735' (Module coreir_or)
  wire [15:0] or_735__in0;
  wire [15:0] or_735__in1;
  wire [15:0] or_735__out;
  coreir_or #(.width(16)) or_735(
    .in0(or_735__in0),
    .in1(or_735__in1),
    .out(or_735__out)
  );

  //Wire declarations for instance 'or_737' (Module coreir_or)
  wire [15:0] or_737__in0;
  wire [15:0] or_737__in1;
  wire [15:0] or_737__out;
  coreir_or #(.width(16)) or_737(
    .in0(or_737__in0),
    .in1(or_737__in1),
    .out(or_737__out)
  );

  //Wire declarations for instance 'or_739' (Module coreir_or)
  wire [15:0] or_739__in0;
  wire [15:0] or_739__in1;
  wire [15:0] or_739__out;
  coreir_or #(.width(16)) or_739(
    .in0(or_739__in0),
    .in1(or_739__in1),
    .out(or_739__out)
  );

  //Wire declarations for instance 'or_741' (Module coreir_or)
  wire [15:0] or_741__in0;
  wire [15:0] or_741__in1;
  wire [15:0] or_741__out;
  coreir_or #(.width(16)) or_741(
    .in0(or_741__in0),
    .in1(or_741__in1),
    .out(or_741__out)
  );

  //Wire declarations for instance 'or_743' (Module coreir_or)
  wire [15:0] or_743__in0;
  wire [15:0] or_743__in1;
  wire [15:0] or_743__out;
  coreir_or #(.width(16)) or_743(
    .in0(or_743__in0),
    .in1(or_743__in1),
    .out(or_743__out)
  );

  //Wire declarations for instance 'or_745' (Module coreir_or)
  wire [15:0] or_745__in0;
  wire [15:0] or_745__in1;
  wire [15:0] or_745__out;
  coreir_or #(.width(16)) or_745(
    .in0(or_745__in0),
    .in1(or_745__in1),
    .out(or_745__out)
  );

  //Wire declarations for instance 'or_747' (Module coreir_or)
  wire [15:0] or_747__in0;
  wire [15:0] or_747__in1;
  wire [15:0] or_747__out;
  coreir_or #(.width(16)) or_747(
    .in0(or_747__in0),
    .in1(or_747__in1),
    .out(or_747__out)
  );

  //Wire declarations for instance 'or_749' (Module coreir_or)
  wire [15:0] or_749__in0;
  wire [15:0] or_749__in1;
  wire [15:0] or_749__out;
  coreir_or #(.width(16)) or_749(
    .in0(or_749__in0),
    .in1(or_749__in1),
    .out(or_749__out)
  );

  //Wire declarations for instance 'or_75' (Module coreir_or)
  wire [15:0] or_75__in0;
  wire [15:0] or_75__in1;
  wire [15:0] or_75__out;
  coreir_or #(.width(16)) or_75(
    .in0(or_75__in0),
    .in1(or_75__in1),
    .out(or_75__out)
  );

  //Wire declarations for instance 'or_751' (Module coreir_or)
  wire [15:0] or_751__in0;
  wire [15:0] or_751__in1;
  wire [15:0] or_751__out;
  coreir_or #(.width(16)) or_751(
    .in0(or_751__in0),
    .in1(or_751__in1),
    .out(or_751__out)
  );

  //Wire declarations for instance 'or_753' (Module coreir_or)
  wire [15:0] or_753__in0;
  wire [15:0] or_753__in1;
  wire [15:0] or_753__out;
  coreir_or #(.width(16)) or_753(
    .in0(or_753__in0),
    .in1(or_753__in1),
    .out(or_753__out)
  );

  //Wire declarations for instance 'or_755' (Module coreir_or)
  wire [15:0] or_755__in0;
  wire [15:0] or_755__in1;
  wire [15:0] or_755__out;
  coreir_or #(.width(16)) or_755(
    .in0(or_755__in0),
    .in1(or_755__in1),
    .out(or_755__out)
  );

  //Wire declarations for instance 'or_757' (Module coreir_or)
  wire [15:0] or_757__in0;
  wire [15:0] or_757__in1;
  wire [15:0] or_757__out;
  coreir_or #(.width(16)) or_757(
    .in0(or_757__in0),
    .in1(or_757__in1),
    .out(or_757__out)
  );

  //Wire declarations for instance 'or_759' (Module coreir_or)
  wire [15:0] or_759__in0;
  wire [15:0] or_759__in1;
  wire [15:0] or_759__out;
  coreir_or #(.width(16)) or_759(
    .in0(or_759__in0),
    .in1(or_759__in1),
    .out(or_759__out)
  );

  //Wire declarations for instance 'or_761' (Module coreir_or)
  wire [15:0] or_761__in0;
  wire [15:0] or_761__in1;
  wire [15:0] or_761__out;
  coreir_or #(.width(16)) or_761(
    .in0(or_761__in0),
    .in1(or_761__in1),
    .out(or_761__out)
  );

  //Wire declarations for instance 'or_763' (Module coreir_or)
  wire [15:0] or_763__in0;
  wire [15:0] or_763__in1;
  wire [15:0] or_763__out;
  coreir_or #(.width(16)) or_763(
    .in0(or_763__in0),
    .in1(or_763__in1),
    .out(or_763__out)
  );

  //Wire declarations for instance 'or_765' (Module coreir_or)
  wire [15:0] or_765__in0;
  wire [15:0] or_765__in1;
  wire [15:0] or_765__out;
  coreir_or #(.width(16)) or_765(
    .in0(or_765__in0),
    .in1(or_765__in1),
    .out(or_765__out)
  );

  //Wire declarations for instance 'or_767' (Module coreir_or)
  wire [15:0] or_767__in0;
  wire [15:0] or_767__in1;
  wire [15:0] or_767__out;
  coreir_or #(.width(16)) or_767(
    .in0(or_767__in0),
    .in1(or_767__in1),
    .out(or_767__out)
  );

  //Wire declarations for instance 'or_769' (Module coreir_or)
  wire [15:0] or_769__in0;
  wire [15:0] or_769__in1;
  wire [15:0] or_769__out;
  coreir_or #(.width(16)) or_769(
    .in0(or_769__in0),
    .in1(or_769__in1),
    .out(or_769__out)
  );

  //Wire declarations for instance 'or_77' (Module coreir_or)
  wire [15:0] or_77__in0;
  wire [15:0] or_77__in1;
  wire [15:0] or_77__out;
  coreir_or #(.width(16)) or_77(
    .in0(or_77__in0),
    .in1(or_77__in1),
    .out(or_77__out)
  );

  //Wire declarations for instance 'or_771' (Module coreir_or)
  wire [15:0] or_771__in0;
  wire [15:0] or_771__in1;
  wire [15:0] or_771__out;
  coreir_or #(.width(16)) or_771(
    .in0(or_771__in0),
    .in1(or_771__in1),
    .out(or_771__out)
  );

  //Wire declarations for instance 'or_773' (Module coreir_or)
  wire [15:0] or_773__in0;
  wire [15:0] or_773__in1;
  wire [15:0] or_773__out;
  coreir_or #(.width(16)) or_773(
    .in0(or_773__in0),
    .in1(or_773__in1),
    .out(or_773__out)
  );

  //Wire declarations for instance 'or_775' (Module coreir_or)
  wire [15:0] or_775__in0;
  wire [15:0] or_775__in1;
  wire [15:0] or_775__out;
  coreir_or #(.width(16)) or_775(
    .in0(or_775__in0),
    .in1(or_775__in1),
    .out(or_775__out)
  );

  //Wire declarations for instance 'or_777' (Module coreir_or)
  wire [15:0] or_777__in0;
  wire [15:0] or_777__in1;
  wire [15:0] or_777__out;
  coreir_or #(.width(16)) or_777(
    .in0(or_777__in0),
    .in1(or_777__in1),
    .out(or_777__out)
  );

  //Wire declarations for instance 'or_779' (Module coreir_or)
  wire [15:0] or_779__in0;
  wire [15:0] or_779__in1;
  wire [15:0] or_779__out;
  coreir_or #(.width(16)) or_779(
    .in0(or_779__in0),
    .in1(or_779__in1),
    .out(or_779__out)
  );

  //Wire declarations for instance 'or_781' (Module coreir_or)
  wire [15:0] or_781__in0;
  wire [15:0] or_781__in1;
  wire [15:0] or_781__out;
  coreir_or #(.width(16)) or_781(
    .in0(or_781__in0),
    .in1(or_781__in1),
    .out(or_781__out)
  );

  //Wire declarations for instance 'or_783' (Module coreir_or)
  wire [15:0] or_783__in0;
  wire [15:0] or_783__in1;
  wire [15:0] or_783__out;
  coreir_or #(.width(16)) or_783(
    .in0(or_783__in0),
    .in1(or_783__in1),
    .out(or_783__out)
  );

  //Wire declarations for instance 'or_785' (Module coreir_or)
  wire [15:0] or_785__in0;
  wire [15:0] or_785__in1;
  wire [15:0] or_785__out;
  coreir_or #(.width(16)) or_785(
    .in0(or_785__in0),
    .in1(or_785__in1),
    .out(or_785__out)
  );

  //Wire declarations for instance 'or_787' (Module coreir_or)
  wire [15:0] or_787__in0;
  wire [15:0] or_787__in1;
  wire [15:0] or_787__out;
  coreir_or #(.width(16)) or_787(
    .in0(or_787__in0),
    .in1(or_787__in1),
    .out(or_787__out)
  );

  //Wire declarations for instance 'or_789' (Module coreir_or)
  wire [15:0] or_789__in0;
  wire [15:0] or_789__in1;
  wire [15:0] or_789__out;
  coreir_or #(.width(16)) or_789(
    .in0(or_789__in0),
    .in1(or_789__in1),
    .out(or_789__out)
  );

  //Wire declarations for instance 'or_79' (Module coreir_or)
  wire [15:0] or_79__in0;
  wire [15:0] or_79__in1;
  wire [15:0] or_79__out;
  coreir_or #(.width(16)) or_79(
    .in0(or_79__in0),
    .in1(or_79__in1),
    .out(or_79__out)
  );

  //Wire declarations for instance 'or_791' (Module coreir_or)
  wire [15:0] or_791__in0;
  wire [15:0] or_791__in1;
  wire [15:0] or_791__out;
  coreir_or #(.width(16)) or_791(
    .in0(or_791__in0),
    .in1(or_791__in1),
    .out(or_791__out)
  );

  //Wire declarations for instance 'or_793' (Module coreir_or)
  wire [15:0] or_793__in0;
  wire [15:0] or_793__in1;
  wire [15:0] or_793__out;
  coreir_or #(.width(16)) or_793(
    .in0(or_793__in0),
    .in1(or_793__in1),
    .out(or_793__out)
  );

  //Wire declarations for instance 'or_795' (Module coreir_or)
  wire [15:0] or_795__in0;
  wire [15:0] or_795__in1;
  wire [15:0] or_795__out;
  coreir_or #(.width(16)) or_795(
    .in0(or_795__in0),
    .in1(or_795__in1),
    .out(or_795__out)
  );

  //Wire declarations for instance 'or_797' (Module coreir_or)
  wire [15:0] or_797__in0;
  wire [15:0] or_797__in1;
  wire [15:0] or_797__out;
  coreir_or #(.width(16)) or_797(
    .in0(or_797__in0),
    .in1(or_797__in1),
    .out(or_797__out)
  );

  //Wire declarations for instance 'or_799' (Module coreir_or)
  wire [15:0] or_799__in0;
  wire [15:0] or_799__in1;
  wire [15:0] or_799__out;
  coreir_or #(.width(16)) or_799(
    .in0(or_799__in0),
    .in1(or_799__in1),
    .out(or_799__out)
  );

  //Wire declarations for instance 'or_801' (Module coreir_or)
  wire [15:0] or_801__in0;
  wire [15:0] or_801__in1;
  wire [15:0] or_801__out;
  coreir_or #(.width(16)) or_801(
    .in0(or_801__in0),
    .in1(or_801__in1),
    .out(or_801__out)
  );

  //Wire declarations for instance 'or_803' (Module coreir_or)
  wire [15:0] or_803__in0;
  wire [15:0] or_803__in1;
  wire [15:0] or_803__out;
  coreir_or #(.width(16)) or_803(
    .in0(or_803__in0),
    .in1(or_803__in1),
    .out(or_803__out)
  );

  //Wire declarations for instance 'or_805' (Module coreir_or)
  wire [15:0] or_805__in0;
  wire [15:0] or_805__in1;
  wire [15:0] or_805__out;
  coreir_or #(.width(16)) or_805(
    .in0(or_805__in0),
    .in1(or_805__in1),
    .out(or_805__out)
  );

  //Wire declarations for instance 'or_807' (Module coreir_or)
  wire [15:0] or_807__in0;
  wire [15:0] or_807__in1;
  wire [15:0] or_807__out;
  coreir_or #(.width(16)) or_807(
    .in0(or_807__in0),
    .in1(or_807__in1),
    .out(or_807__out)
  );

  //Wire declarations for instance 'or_809' (Module coreir_or)
  wire [15:0] or_809__in0;
  wire [15:0] or_809__in1;
  wire [15:0] or_809__out;
  coreir_or #(.width(16)) or_809(
    .in0(or_809__in0),
    .in1(or_809__in1),
    .out(or_809__out)
  );

  //Wire declarations for instance 'or_81' (Module coreir_or)
  wire [15:0] or_81__in0;
  wire [15:0] or_81__in1;
  wire [15:0] or_81__out;
  coreir_or #(.width(16)) or_81(
    .in0(or_81__in0),
    .in1(or_81__in1),
    .out(or_81__out)
  );

  //Wire declarations for instance 'or_811' (Module coreir_or)
  wire [15:0] or_811__in0;
  wire [15:0] or_811__in1;
  wire [15:0] or_811__out;
  coreir_or #(.width(16)) or_811(
    .in0(or_811__in0),
    .in1(or_811__in1),
    .out(or_811__out)
  );

  //Wire declarations for instance 'or_813' (Module coreir_or)
  wire [15:0] or_813__in0;
  wire [15:0] or_813__in1;
  wire [15:0] or_813__out;
  coreir_or #(.width(16)) or_813(
    .in0(or_813__in0),
    .in1(or_813__in1),
    .out(or_813__out)
  );

  //Wire declarations for instance 'or_815' (Module coreir_or)
  wire [15:0] or_815__in0;
  wire [15:0] or_815__in1;
  wire [15:0] or_815__out;
  coreir_or #(.width(16)) or_815(
    .in0(or_815__in0),
    .in1(or_815__in1),
    .out(or_815__out)
  );

  //Wire declarations for instance 'or_817' (Module coreir_or)
  wire [15:0] or_817__in0;
  wire [15:0] or_817__in1;
  wire [15:0] or_817__out;
  coreir_or #(.width(16)) or_817(
    .in0(or_817__in0),
    .in1(or_817__in1),
    .out(or_817__out)
  );

  //Wire declarations for instance 'or_819' (Module coreir_or)
  wire [15:0] or_819__in0;
  wire [15:0] or_819__in1;
  wire [15:0] or_819__out;
  coreir_or #(.width(16)) or_819(
    .in0(or_819__in0),
    .in1(or_819__in1),
    .out(or_819__out)
  );

  //Wire declarations for instance 'or_821' (Module coreir_or)
  wire [15:0] or_821__in0;
  wire [15:0] or_821__in1;
  wire [15:0] or_821__out;
  coreir_or #(.width(16)) or_821(
    .in0(or_821__in0),
    .in1(or_821__in1),
    .out(or_821__out)
  );

  //Wire declarations for instance 'or_823' (Module coreir_or)
  wire [15:0] or_823__in0;
  wire [15:0] or_823__in1;
  wire [15:0] or_823__out;
  coreir_or #(.width(16)) or_823(
    .in0(or_823__in0),
    .in1(or_823__in1),
    .out(or_823__out)
  );

  //Wire declarations for instance 'or_825' (Module coreir_or)
  wire [15:0] or_825__in0;
  wire [15:0] or_825__in1;
  wire [15:0] or_825__out;
  coreir_or #(.width(16)) or_825(
    .in0(or_825__in0),
    .in1(or_825__in1),
    .out(or_825__out)
  );

  //Wire declarations for instance 'or_827' (Module coreir_or)
  wire [15:0] or_827__in0;
  wire [15:0] or_827__in1;
  wire [15:0] or_827__out;
  coreir_or #(.width(16)) or_827(
    .in0(or_827__in0),
    .in1(or_827__in1),
    .out(or_827__out)
  );

  //Wire declarations for instance 'or_829' (Module coreir_or)
  wire [15:0] or_829__in0;
  wire [15:0] or_829__in1;
  wire [15:0] or_829__out;
  coreir_or #(.width(16)) or_829(
    .in0(or_829__in0),
    .in1(or_829__in1),
    .out(or_829__out)
  );

  //Wire declarations for instance 'or_83' (Module coreir_or)
  wire [15:0] or_83__in0;
  wire [15:0] or_83__in1;
  wire [15:0] or_83__out;
  coreir_or #(.width(16)) or_83(
    .in0(or_83__in0),
    .in1(or_83__in1),
    .out(or_83__out)
  );

  //Wire declarations for instance 'or_831' (Module coreir_or)
  wire [15:0] or_831__in0;
  wire [15:0] or_831__in1;
  wire [15:0] or_831__out;
  coreir_or #(.width(16)) or_831(
    .in0(or_831__in0),
    .in1(or_831__in1),
    .out(or_831__out)
  );

  //Wire declarations for instance 'or_833' (Module coreir_or)
  wire [15:0] or_833__in0;
  wire [15:0] or_833__in1;
  wire [15:0] or_833__out;
  coreir_or #(.width(16)) or_833(
    .in0(or_833__in0),
    .in1(or_833__in1),
    .out(or_833__out)
  );

  //Wire declarations for instance 'or_835' (Module coreir_or)
  wire [15:0] or_835__in0;
  wire [15:0] or_835__in1;
  wire [15:0] or_835__out;
  coreir_or #(.width(16)) or_835(
    .in0(or_835__in0),
    .in1(or_835__in1),
    .out(or_835__out)
  );

  //Wire declarations for instance 'or_837' (Module coreir_or)
  wire [15:0] or_837__in0;
  wire [15:0] or_837__in1;
  wire [15:0] or_837__out;
  coreir_or #(.width(16)) or_837(
    .in0(or_837__in0),
    .in1(or_837__in1),
    .out(or_837__out)
  );

  //Wire declarations for instance 'or_839' (Module coreir_or)
  wire [15:0] or_839__in0;
  wire [15:0] or_839__in1;
  wire [15:0] or_839__out;
  coreir_or #(.width(16)) or_839(
    .in0(or_839__in0),
    .in1(or_839__in1),
    .out(or_839__out)
  );

  //Wire declarations for instance 'or_841' (Module coreir_or)
  wire [15:0] or_841__in0;
  wire [15:0] or_841__in1;
  wire [15:0] or_841__out;
  coreir_or #(.width(16)) or_841(
    .in0(or_841__in0),
    .in1(or_841__in1),
    .out(or_841__out)
  );

  //Wire declarations for instance 'or_843' (Module coreir_or)
  wire [15:0] or_843__in0;
  wire [15:0] or_843__in1;
  wire [15:0] or_843__out;
  coreir_or #(.width(16)) or_843(
    .in0(or_843__in0),
    .in1(or_843__in1),
    .out(or_843__out)
  );

  //Wire declarations for instance 'or_845' (Module coreir_or)
  wire [15:0] or_845__in0;
  wire [15:0] or_845__in1;
  wire [15:0] or_845__out;
  coreir_or #(.width(16)) or_845(
    .in0(or_845__in0),
    .in1(or_845__in1),
    .out(or_845__out)
  );

  //Wire declarations for instance 'or_847' (Module coreir_or)
  wire [15:0] or_847__in0;
  wire [15:0] or_847__in1;
  wire [15:0] or_847__out;
  coreir_or #(.width(16)) or_847(
    .in0(or_847__in0),
    .in1(or_847__in1),
    .out(or_847__out)
  );

  //Wire declarations for instance 'or_849' (Module coreir_or)
  wire [15:0] or_849__in0;
  wire [15:0] or_849__in1;
  wire [15:0] or_849__out;
  coreir_or #(.width(16)) or_849(
    .in0(or_849__in0),
    .in1(or_849__in1),
    .out(or_849__out)
  );

  //Wire declarations for instance 'or_85' (Module coreir_or)
  wire [15:0] or_85__in0;
  wire [15:0] or_85__in1;
  wire [15:0] or_85__out;
  coreir_or #(.width(16)) or_85(
    .in0(or_85__in0),
    .in1(or_85__in1),
    .out(or_85__out)
  );

  //Wire declarations for instance 'or_851' (Module coreir_or)
  wire [15:0] or_851__in0;
  wire [15:0] or_851__in1;
  wire [15:0] or_851__out;
  coreir_or #(.width(16)) or_851(
    .in0(or_851__in0),
    .in1(or_851__in1),
    .out(or_851__out)
  );

  //Wire declarations for instance 'or_853' (Module coreir_or)
  wire [15:0] or_853__in0;
  wire [15:0] or_853__in1;
  wire [15:0] or_853__out;
  coreir_or #(.width(16)) or_853(
    .in0(or_853__in0),
    .in1(or_853__in1),
    .out(or_853__out)
  );

  //Wire declarations for instance 'or_855' (Module coreir_or)
  wire [15:0] or_855__in0;
  wire [15:0] or_855__in1;
  wire [15:0] or_855__out;
  coreir_or #(.width(16)) or_855(
    .in0(or_855__in0),
    .in1(or_855__in1),
    .out(or_855__out)
  );

  //Wire declarations for instance 'or_857' (Module coreir_or)
  wire [15:0] or_857__in0;
  wire [15:0] or_857__in1;
  wire [15:0] or_857__out;
  coreir_or #(.width(16)) or_857(
    .in0(or_857__in0),
    .in1(or_857__in1),
    .out(or_857__out)
  );

  //Wire declarations for instance 'or_859' (Module coreir_or)
  wire [15:0] or_859__in0;
  wire [15:0] or_859__in1;
  wire [15:0] or_859__out;
  coreir_or #(.width(16)) or_859(
    .in0(or_859__in0),
    .in1(or_859__in1),
    .out(or_859__out)
  );

  //Wire declarations for instance 'or_861' (Module coreir_or)
  wire [15:0] or_861__in0;
  wire [15:0] or_861__in1;
  wire [15:0] or_861__out;
  coreir_or #(.width(16)) or_861(
    .in0(or_861__in0),
    .in1(or_861__in1),
    .out(or_861__out)
  );

  //Wire declarations for instance 'or_863' (Module coreir_or)
  wire [15:0] or_863__in0;
  wire [15:0] or_863__in1;
  wire [15:0] or_863__out;
  coreir_or #(.width(16)) or_863(
    .in0(or_863__in0),
    .in1(or_863__in1),
    .out(or_863__out)
  );

  //Wire declarations for instance 'or_865' (Module coreir_or)
  wire [15:0] or_865__in0;
  wire [15:0] or_865__in1;
  wire [15:0] or_865__out;
  coreir_or #(.width(16)) or_865(
    .in0(or_865__in0),
    .in1(or_865__in1),
    .out(or_865__out)
  );

  //Wire declarations for instance 'or_867' (Module coreir_or)
  wire [15:0] or_867__in0;
  wire [15:0] or_867__in1;
  wire [15:0] or_867__out;
  coreir_or #(.width(16)) or_867(
    .in0(or_867__in0),
    .in1(or_867__in1),
    .out(or_867__out)
  );

  //Wire declarations for instance 'or_869' (Module coreir_or)
  wire [15:0] or_869__in0;
  wire [15:0] or_869__in1;
  wire [15:0] or_869__out;
  coreir_or #(.width(16)) or_869(
    .in0(or_869__in0),
    .in1(or_869__in1),
    .out(or_869__out)
  );

  //Wire declarations for instance 'or_87' (Module coreir_or)
  wire [15:0] or_87__in0;
  wire [15:0] or_87__in1;
  wire [15:0] or_87__out;
  coreir_or #(.width(16)) or_87(
    .in0(or_87__in0),
    .in1(or_87__in1),
    .out(or_87__out)
  );

  //Wire declarations for instance 'or_871' (Module coreir_or)
  wire [15:0] or_871__in0;
  wire [15:0] or_871__in1;
  wire [15:0] or_871__out;
  coreir_or #(.width(16)) or_871(
    .in0(or_871__in0),
    .in1(or_871__in1),
    .out(or_871__out)
  );

  //Wire declarations for instance 'or_873' (Module coreir_or)
  wire [15:0] or_873__in0;
  wire [15:0] or_873__in1;
  wire [15:0] or_873__out;
  coreir_or #(.width(16)) or_873(
    .in0(or_873__in0),
    .in1(or_873__in1),
    .out(or_873__out)
  );

  //Wire declarations for instance 'or_875' (Module coreir_or)
  wire [15:0] or_875__in0;
  wire [15:0] or_875__in1;
  wire [15:0] or_875__out;
  coreir_or #(.width(16)) or_875(
    .in0(or_875__in0),
    .in1(or_875__in1),
    .out(or_875__out)
  );

  //Wire declarations for instance 'or_877' (Module coreir_or)
  wire [15:0] or_877__in0;
  wire [15:0] or_877__in1;
  wire [15:0] or_877__out;
  coreir_or #(.width(16)) or_877(
    .in0(or_877__in0),
    .in1(or_877__in1),
    .out(or_877__out)
  );

  //Wire declarations for instance 'or_879' (Module coreir_or)
  wire [15:0] or_879__in0;
  wire [15:0] or_879__in1;
  wire [15:0] or_879__out;
  coreir_or #(.width(16)) or_879(
    .in0(or_879__in0),
    .in1(or_879__in1),
    .out(or_879__out)
  );

  //Wire declarations for instance 'or_881' (Module coreir_or)
  wire [15:0] or_881__in0;
  wire [15:0] or_881__in1;
  wire [15:0] or_881__out;
  coreir_or #(.width(16)) or_881(
    .in0(or_881__in0),
    .in1(or_881__in1),
    .out(or_881__out)
  );

  //Wire declarations for instance 'or_883' (Module coreir_or)
  wire [15:0] or_883__in0;
  wire [15:0] or_883__in1;
  wire [15:0] or_883__out;
  coreir_or #(.width(16)) or_883(
    .in0(or_883__in0),
    .in1(or_883__in1),
    .out(or_883__out)
  );

  //Wire declarations for instance 'or_885' (Module coreir_or)
  wire [15:0] or_885__in0;
  wire [15:0] or_885__in1;
  wire [15:0] or_885__out;
  coreir_or #(.width(16)) or_885(
    .in0(or_885__in0),
    .in1(or_885__in1),
    .out(or_885__out)
  );

  //Wire declarations for instance 'or_887' (Module coreir_or)
  wire [15:0] or_887__in0;
  wire [15:0] or_887__in1;
  wire [15:0] or_887__out;
  coreir_or #(.width(16)) or_887(
    .in0(or_887__in0),
    .in1(or_887__in1),
    .out(or_887__out)
  );

  //Wire declarations for instance 'or_889' (Module coreir_or)
  wire [15:0] or_889__in0;
  wire [15:0] or_889__in1;
  wire [15:0] or_889__out;
  coreir_or #(.width(16)) or_889(
    .in0(or_889__in0),
    .in1(or_889__in1),
    .out(or_889__out)
  );

  //Wire declarations for instance 'or_89' (Module coreir_or)
  wire [15:0] or_89__in0;
  wire [15:0] or_89__in1;
  wire [15:0] or_89__out;
  coreir_or #(.width(16)) or_89(
    .in0(or_89__in0),
    .in1(or_89__in1),
    .out(or_89__out)
  );

  //Wire declarations for instance 'or_891' (Module coreir_or)
  wire [15:0] or_891__in0;
  wire [15:0] or_891__in1;
  wire [15:0] or_891__out;
  coreir_or #(.width(16)) or_891(
    .in0(or_891__in0),
    .in1(or_891__in1),
    .out(or_891__out)
  );

  //Wire declarations for instance 'or_893' (Module coreir_or)
  wire [15:0] or_893__in0;
  wire [15:0] or_893__in1;
  wire [15:0] or_893__out;
  coreir_or #(.width(16)) or_893(
    .in0(or_893__in0),
    .in1(or_893__in1),
    .out(or_893__out)
  );

  //Wire declarations for instance 'or_895' (Module coreir_or)
  wire [15:0] or_895__in0;
  wire [15:0] or_895__in1;
  wire [15:0] or_895__out;
  coreir_or #(.width(16)) or_895(
    .in0(or_895__in0),
    .in1(or_895__in1),
    .out(or_895__out)
  );

  //Wire declarations for instance 'or_897' (Module coreir_or)
  wire [15:0] or_897__in0;
  wire [15:0] or_897__in1;
  wire [15:0] or_897__out;
  coreir_or #(.width(16)) or_897(
    .in0(or_897__in0),
    .in1(or_897__in1),
    .out(or_897__out)
  );

  //Wire declarations for instance 'or_899' (Module coreir_or)
  wire [15:0] or_899__in0;
  wire [15:0] or_899__in1;
  wire [15:0] or_899__out;
  coreir_or #(.width(16)) or_899(
    .in0(or_899__in0),
    .in1(or_899__in1),
    .out(or_899__out)
  );

  //Wire declarations for instance 'or_9' (Module coreir_or)
  wire [15:0] or_9__in0;
  wire [15:0] or_9__in1;
  wire [15:0] or_9__out;
  coreir_or #(.width(16)) or_9(
    .in0(or_9__in0),
    .in1(or_9__in1),
    .out(or_9__out)
  );

  //Wire declarations for instance 'or_901' (Module coreir_or)
  wire [15:0] or_901__in0;
  wire [15:0] or_901__in1;
  wire [15:0] or_901__out;
  coreir_or #(.width(16)) or_901(
    .in0(or_901__in0),
    .in1(or_901__in1),
    .out(or_901__out)
  );

  //Wire declarations for instance 'or_903' (Module coreir_or)
  wire [15:0] or_903__in0;
  wire [15:0] or_903__in1;
  wire [15:0] or_903__out;
  coreir_or #(.width(16)) or_903(
    .in0(or_903__in0),
    .in1(or_903__in1),
    .out(or_903__out)
  );

  //Wire declarations for instance 'or_905' (Module coreir_or)
  wire [15:0] or_905__in0;
  wire [15:0] or_905__in1;
  wire [15:0] or_905__out;
  coreir_or #(.width(16)) or_905(
    .in0(or_905__in0),
    .in1(or_905__in1),
    .out(or_905__out)
  );

  //Wire declarations for instance 'or_907' (Module coreir_or)
  wire [15:0] or_907__in0;
  wire [15:0] or_907__in1;
  wire [15:0] or_907__out;
  coreir_or #(.width(16)) or_907(
    .in0(or_907__in0),
    .in1(or_907__in1),
    .out(or_907__out)
  );

  //Wire declarations for instance 'or_909' (Module coreir_or)
  wire [15:0] or_909__in0;
  wire [15:0] or_909__in1;
  wire [15:0] or_909__out;
  coreir_or #(.width(16)) or_909(
    .in0(or_909__in0),
    .in1(or_909__in1),
    .out(or_909__out)
  );

  //Wire declarations for instance 'or_91' (Module coreir_or)
  wire [15:0] or_91__in0;
  wire [15:0] or_91__in1;
  wire [15:0] or_91__out;
  coreir_or #(.width(16)) or_91(
    .in0(or_91__in0),
    .in1(or_91__in1),
    .out(or_91__out)
  );

  //Wire declarations for instance 'or_911' (Module coreir_or)
  wire [15:0] or_911__in0;
  wire [15:0] or_911__in1;
  wire [15:0] or_911__out;
  coreir_or #(.width(16)) or_911(
    .in0(or_911__in0),
    .in1(or_911__in1),
    .out(or_911__out)
  );

  //Wire declarations for instance 'or_913' (Module coreir_or)
  wire [15:0] or_913__in0;
  wire [15:0] or_913__in1;
  wire [15:0] or_913__out;
  coreir_or #(.width(16)) or_913(
    .in0(or_913__in0),
    .in1(or_913__in1),
    .out(or_913__out)
  );

  //Wire declarations for instance 'or_915' (Module coreir_or)
  wire [15:0] or_915__in0;
  wire [15:0] or_915__in1;
  wire [15:0] or_915__out;
  coreir_or #(.width(16)) or_915(
    .in0(or_915__in0),
    .in1(or_915__in1),
    .out(or_915__out)
  );

  //Wire declarations for instance 'or_917' (Module coreir_or)
  wire [15:0] or_917__in0;
  wire [15:0] or_917__in1;
  wire [15:0] or_917__out;
  coreir_or #(.width(16)) or_917(
    .in0(or_917__in0),
    .in1(or_917__in1),
    .out(or_917__out)
  );

  //Wire declarations for instance 'or_919' (Module coreir_or)
  wire [15:0] or_919__in0;
  wire [15:0] or_919__in1;
  wire [15:0] or_919__out;
  coreir_or #(.width(16)) or_919(
    .in0(or_919__in0),
    .in1(or_919__in1),
    .out(or_919__out)
  );

  //Wire declarations for instance 'or_921' (Module coreir_or)
  wire [15:0] or_921__in0;
  wire [15:0] or_921__in1;
  wire [15:0] or_921__out;
  coreir_or #(.width(16)) or_921(
    .in0(or_921__in0),
    .in1(or_921__in1),
    .out(or_921__out)
  );

  //Wire declarations for instance 'or_923' (Module coreir_or)
  wire [15:0] or_923__in0;
  wire [15:0] or_923__in1;
  wire [15:0] or_923__out;
  coreir_or #(.width(16)) or_923(
    .in0(or_923__in0),
    .in1(or_923__in1),
    .out(or_923__out)
  );

  //Wire declarations for instance 'or_925' (Module coreir_or)
  wire [15:0] or_925__in0;
  wire [15:0] or_925__in1;
  wire [15:0] or_925__out;
  coreir_or #(.width(16)) or_925(
    .in0(or_925__in0),
    .in1(or_925__in1),
    .out(or_925__out)
  );

  //Wire declarations for instance 'or_927' (Module coreir_or)
  wire [15:0] or_927__in0;
  wire [15:0] or_927__in1;
  wire [15:0] or_927__out;
  coreir_or #(.width(16)) or_927(
    .in0(or_927__in0),
    .in1(or_927__in1),
    .out(or_927__out)
  );

  //Wire declarations for instance 'or_929' (Module coreir_or)
  wire [15:0] or_929__in0;
  wire [15:0] or_929__in1;
  wire [15:0] or_929__out;
  coreir_or #(.width(16)) or_929(
    .in0(or_929__in0),
    .in1(or_929__in1),
    .out(or_929__out)
  );

  //Wire declarations for instance 'or_93' (Module coreir_or)
  wire [15:0] or_93__in0;
  wire [15:0] or_93__in1;
  wire [15:0] or_93__out;
  coreir_or #(.width(16)) or_93(
    .in0(or_93__in0),
    .in1(or_93__in1),
    .out(or_93__out)
  );

  //Wire declarations for instance 'or_931' (Module coreir_or)
  wire [15:0] or_931__in0;
  wire [15:0] or_931__in1;
  wire [15:0] or_931__out;
  coreir_or #(.width(16)) or_931(
    .in0(or_931__in0),
    .in1(or_931__in1),
    .out(or_931__out)
  );

  //Wire declarations for instance 'or_933' (Module coreir_or)
  wire [15:0] or_933__in0;
  wire [15:0] or_933__in1;
  wire [15:0] or_933__out;
  coreir_or #(.width(16)) or_933(
    .in0(or_933__in0),
    .in1(or_933__in1),
    .out(or_933__out)
  );

  //Wire declarations for instance 'or_935' (Module coreir_or)
  wire [15:0] or_935__in0;
  wire [15:0] or_935__in1;
  wire [15:0] or_935__out;
  coreir_or #(.width(16)) or_935(
    .in0(or_935__in0),
    .in1(or_935__in1),
    .out(or_935__out)
  );

  //Wire declarations for instance 'or_937' (Module coreir_or)
  wire [15:0] or_937__in0;
  wire [15:0] or_937__in1;
  wire [15:0] or_937__out;
  coreir_or #(.width(16)) or_937(
    .in0(or_937__in0),
    .in1(or_937__in1),
    .out(or_937__out)
  );

  //Wire declarations for instance 'or_939' (Module coreir_or)
  wire [15:0] or_939__in0;
  wire [15:0] or_939__in1;
  wire [15:0] or_939__out;
  coreir_or #(.width(16)) or_939(
    .in0(or_939__in0),
    .in1(or_939__in1),
    .out(or_939__out)
  );

  //Wire declarations for instance 'or_941' (Module coreir_or)
  wire [15:0] or_941__in0;
  wire [15:0] or_941__in1;
  wire [15:0] or_941__out;
  coreir_or #(.width(16)) or_941(
    .in0(or_941__in0),
    .in1(or_941__in1),
    .out(or_941__out)
  );

  //Wire declarations for instance 'or_943' (Module coreir_or)
  wire [15:0] or_943__in0;
  wire [15:0] or_943__in1;
  wire [15:0] or_943__out;
  coreir_or #(.width(16)) or_943(
    .in0(or_943__in0),
    .in1(or_943__in1),
    .out(or_943__out)
  );

  //Wire declarations for instance 'or_945' (Module coreir_or)
  wire [15:0] or_945__in0;
  wire [15:0] or_945__in1;
  wire [15:0] or_945__out;
  coreir_or #(.width(16)) or_945(
    .in0(or_945__in0),
    .in1(or_945__in1),
    .out(or_945__out)
  );

  //Wire declarations for instance 'or_947' (Module coreir_or)
  wire [15:0] or_947__in0;
  wire [15:0] or_947__in1;
  wire [15:0] or_947__out;
  coreir_or #(.width(16)) or_947(
    .in0(or_947__in0),
    .in1(or_947__in1),
    .out(or_947__out)
  );

  //Wire declarations for instance 'or_949' (Module coreir_or)
  wire [15:0] or_949__in0;
  wire [15:0] or_949__in1;
  wire [15:0] or_949__out;
  coreir_or #(.width(16)) or_949(
    .in0(or_949__in0),
    .in1(or_949__in1),
    .out(or_949__out)
  );

  //Wire declarations for instance 'or_95' (Module coreir_or)
  wire [15:0] or_95__in0;
  wire [15:0] or_95__in1;
  wire [15:0] or_95__out;
  coreir_or #(.width(16)) or_95(
    .in0(or_95__in0),
    .in1(or_95__in1),
    .out(or_95__out)
  );

  //Wire declarations for instance 'or_951' (Module coreir_or)
  wire [15:0] or_951__in0;
  wire [15:0] or_951__in1;
  wire [15:0] or_951__out;
  coreir_or #(.width(16)) or_951(
    .in0(or_951__in0),
    .in1(or_951__in1),
    .out(or_951__out)
  );

  //Wire declarations for instance 'or_953' (Module coreir_or)
  wire [15:0] or_953__in0;
  wire [15:0] or_953__in1;
  wire [15:0] or_953__out;
  coreir_or #(.width(16)) or_953(
    .in0(or_953__in0),
    .in1(or_953__in1),
    .out(or_953__out)
  );

  //Wire declarations for instance 'or_955' (Module coreir_or)
  wire [15:0] or_955__in0;
  wire [15:0] or_955__in1;
  wire [15:0] or_955__out;
  coreir_or #(.width(16)) or_955(
    .in0(or_955__in0),
    .in1(or_955__in1),
    .out(or_955__out)
  );

  //Wire declarations for instance 'or_957' (Module coreir_or)
  wire [15:0] or_957__in0;
  wire [15:0] or_957__in1;
  wire [15:0] or_957__out;
  coreir_or #(.width(16)) or_957(
    .in0(or_957__in0),
    .in1(or_957__in1),
    .out(or_957__out)
  );

  //Wire declarations for instance 'or_959' (Module coreir_or)
  wire [15:0] or_959__in0;
  wire [15:0] or_959__in1;
  wire [15:0] or_959__out;
  coreir_or #(.width(16)) or_959(
    .in0(or_959__in0),
    .in1(or_959__in1),
    .out(or_959__out)
  );

  //Wire declarations for instance 'or_961' (Module coreir_or)
  wire [15:0] or_961__in0;
  wire [15:0] or_961__in1;
  wire [15:0] or_961__out;
  coreir_or #(.width(16)) or_961(
    .in0(or_961__in0),
    .in1(or_961__in1),
    .out(or_961__out)
  );

  //Wire declarations for instance 'or_963' (Module coreir_or)
  wire [15:0] or_963__in0;
  wire [15:0] or_963__in1;
  wire [15:0] or_963__out;
  coreir_or #(.width(16)) or_963(
    .in0(or_963__in0),
    .in1(or_963__in1),
    .out(or_963__out)
  );

  //Wire declarations for instance 'or_965' (Module coreir_or)
  wire [15:0] or_965__in0;
  wire [15:0] or_965__in1;
  wire [15:0] or_965__out;
  coreir_or #(.width(16)) or_965(
    .in0(or_965__in0),
    .in1(or_965__in1),
    .out(or_965__out)
  );

  //Wire declarations for instance 'or_967' (Module coreir_or)
  wire [15:0] or_967__in0;
  wire [15:0] or_967__in1;
  wire [15:0] or_967__out;
  coreir_or #(.width(16)) or_967(
    .in0(or_967__in0),
    .in1(or_967__in1),
    .out(or_967__out)
  );

  //Wire declarations for instance 'or_969' (Module coreir_or)
  wire [15:0] or_969__in0;
  wire [15:0] or_969__in1;
  wire [15:0] or_969__out;
  coreir_or #(.width(16)) or_969(
    .in0(or_969__in0),
    .in1(or_969__in1),
    .out(or_969__out)
  );

  //Wire declarations for instance 'or_97' (Module coreir_or)
  wire [15:0] or_97__in0;
  wire [15:0] or_97__in1;
  wire [15:0] or_97__out;
  coreir_or #(.width(16)) or_97(
    .in0(or_97__in0),
    .in1(or_97__in1),
    .out(or_97__out)
  );

  //Wire declarations for instance 'or_971' (Module coreir_or)
  wire [15:0] or_971__in0;
  wire [15:0] or_971__in1;
  wire [15:0] or_971__out;
  coreir_or #(.width(16)) or_971(
    .in0(or_971__in0),
    .in1(or_971__in1),
    .out(or_971__out)
  );

  //Wire declarations for instance 'or_973' (Module coreir_or)
  wire [15:0] or_973__in0;
  wire [15:0] or_973__in1;
  wire [15:0] or_973__out;
  coreir_or #(.width(16)) or_973(
    .in0(or_973__in0),
    .in1(or_973__in1),
    .out(or_973__out)
  );

  //Wire declarations for instance 'or_975' (Module coreir_or)
  wire [15:0] or_975__in0;
  wire [15:0] or_975__in1;
  wire [15:0] or_975__out;
  coreir_or #(.width(16)) or_975(
    .in0(or_975__in0),
    .in1(or_975__in1),
    .out(or_975__out)
  );

  //Wire declarations for instance 'or_977' (Module coreir_or)
  wire [15:0] or_977__in0;
  wire [15:0] or_977__in1;
  wire [15:0] or_977__out;
  coreir_or #(.width(16)) or_977(
    .in0(or_977__in0),
    .in1(or_977__in1),
    .out(or_977__out)
  );

  //Wire declarations for instance 'or_979' (Module coreir_or)
  wire [15:0] or_979__in0;
  wire [15:0] or_979__in1;
  wire [15:0] or_979__out;
  coreir_or #(.width(16)) or_979(
    .in0(or_979__in0),
    .in1(or_979__in1),
    .out(or_979__out)
  );

  //Wire declarations for instance 'or_981' (Module coreir_or)
  wire [15:0] or_981__in0;
  wire [15:0] or_981__in1;
  wire [15:0] or_981__out;
  coreir_or #(.width(16)) or_981(
    .in0(or_981__in0),
    .in1(or_981__in1),
    .out(or_981__out)
  );

  //Wire declarations for instance 'or_983' (Module coreir_or)
  wire [15:0] or_983__in0;
  wire [15:0] or_983__in1;
  wire [15:0] or_983__out;
  coreir_or #(.width(16)) or_983(
    .in0(or_983__in0),
    .in1(or_983__in1),
    .out(or_983__out)
  );

  //Wire declarations for instance 'or_985' (Module coreir_or)
  wire [15:0] or_985__in0;
  wire [15:0] or_985__in1;
  wire [15:0] or_985__out;
  coreir_or #(.width(16)) or_985(
    .in0(or_985__in0),
    .in1(or_985__in1),
    .out(or_985__out)
  );

  //Wire declarations for instance 'or_987' (Module coreir_or)
  wire [15:0] or_987__in0;
  wire [15:0] or_987__in1;
  wire [15:0] or_987__out;
  coreir_or #(.width(16)) or_987(
    .in0(or_987__in0),
    .in1(or_987__in1),
    .out(or_987__out)
  );

  //Wire declarations for instance 'or_989' (Module coreir_or)
  wire [15:0] or_989__in0;
  wire [15:0] or_989__in1;
  wire [15:0] or_989__out;
  coreir_or #(.width(16)) or_989(
    .in0(or_989__in0),
    .in1(or_989__in1),
    .out(or_989__out)
  );

  //Wire declarations for instance 'or_99' (Module coreir_or)
  wire [15:0] or_99__in0;
  wire [15:0] or_99__in1;
  wire [15:0] or_99__out;
  coreir_or #(.width(16)) or_99(
    .in0(or_99__in0),
    .in1(or_99__in1),
    .out(or_99__out)
  );

  //Wire declarations for instance 'or_991' (Module coreir_or)
  wire [15:0] or_991__in0;
  wire [15:0] or_991__in1;
  wire [15:0] or_991__out;
  coreir_or #(.width(16)) or_991(
    .in0(or_991__in0),
    .in1(or_991__in1),
    .out(or_991__out)
  );

  //Wire declarations for instance 'or_993' (Module coreir_or)
  wire [15:0] or_993__in0;
  wire [15:0] or_993__in1;
  wire [15:0] or_993__out;
  coreir_or #(.width(16)) or_993(
    .in0(or_993__in0),
    .in1(or_993__in1),
    .out(or_993__out)
  );

  //Wire declarations for instance 'or_995' (Module coreir_or)
  wire [15:0] or_995__in0;
  wire [15:0] or_995__in1;
  wire [15:0] or_995__out;
  coreir_or #(.width(16)) or_995(
    .in0(or_995__in0),
    .in1(or_995__in1),
    .out(or_995__out)
  );

  //Wire declarations for instance 'or_997' (Module coreir_or)
  wire [15:0] or_997__in0;
  wire [15:0] or_997__in1;
  wire [15:0] or_997__out;
  coreir_or #(.width(16)) or_997(
    .in0(or_997__in0),
    .in1(or_997__in1),
    .out(or_997__out)
  );

  //Wire declarations for instance 'or_999' (Module coreir_or)
  wire [15:0] or_999__in0;
  wire [15:0] or_999__in1;
  wire [15:0] or_999__out;
  coreir_or #(.width(16)) or_999(
    .in0(or_999__in0),
    .in1(or_999__in1),
    .out(or_999__out)
  );

  //Wire declarations for instance 'reg_0' (Module coreir_reg)
  wire  reg_0__clk;
  wire [15:0] reg_0__in;
  wire [15:0] reg_0__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_0(
    .clk(reg_0__clk),
    .in(reg_0__in),
    .out(reg_0__out)
  );

  //Wire declarations for instance 'reg_1' (Module coreir_reg)
  wire  reg_1__clk;
  wire [15:0] reg_1__in;
  wire [15:0] reg_1__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_1(
    .clk(reg_1__clk),
    .in(reg_1__in),
    .out(reg_1__out)
  );

  //Wire declarations for instance 'reg_10' (Module coreir_reg)
  wire  reg_10__clk;
  wire [15:0] reg_10__in;
  wire [15:0] reg_10__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_10(
    .clk(reg_10__clk),
    .in(reg_10__in),
    .out(reg_10__out)
  );

  //Wire declarations for instance 'reg_100' (Module coreir_reg)
  wire  reg_100__clk;
  wire [15:0] reg_100__in;
  wire [15:0] reg_100__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_100(
    .clk(reg_100__clk),
    .in(reg_100__in),
    .out(reg_100__out)
  );

  //Wire declarations for instance 'reg_101' (Module coreir_reg)
  wire  reg_101__clk;
  wire [15:0] reg_101__in;
  wire [15:0] reg_101__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_101(
    .clk(reg_101__clk),
    .in(reg_101__in),
    .out(reg_101__out)
  );

  //Wire declarations for instance 'reg_102' (Module coreir_reg)
  wire  reg_102__clk;
  wire [15:0] reg_102__in;
  wire [15:0] reg_102__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_102(
    .clk(reg_102__clk),
    .in(reg_102__in),
    .out(reg_102__out)
  );

  //Wire declarations for instance 'reg_103' (Module coreir_reg)
  wire  reg_103__clk;
  wire [15:0] reg_103__in;
  wire [15:0] reg_103__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_103(
    .clk(reg_103__clk),
    .in(reg_103__in),
    .out(reg_103__out)
  );

  //Wire declarations for instance 'reg_104' (Module coreir_reg)
  wire  reg_104__clk;
  wire [15:0] reg_104__in;
  wire [15:0] reg_104__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_104(
    .clk(reg_104__clk),
    .in(reg_104__in),
    .out(reg_104__out)
  );

  //Wire declarations for instance 'reg_105' (Module coreir_reg)
  wire  reg_105__clk;
  wire [15:0] reg_105__in;
  wire [15:0] reg_105__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_105(
    .clk(reg_105__clk),
    .in(reg_105__in),
    .out(reg_105__out)
  );

  //Wire declarations for instance 'reg_106' (Module coreir_reg)
  wire  reg_106__clk;
  wire [15:0] reg_106__in;
  wire [15:0] reg_106__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_106(
    .clk(reg_106__clk),
    .in(reg_106__in),
    .out(reg_106__out)
  );

  //Wire declarations for instance 'reg_107' (Module coreir_reg)
  wire  reg_107__clk;
  wire [15:0] reg_107__in;
  wire [15:0] reg_107__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_107(
    .clk(reg_107__clk),
    .in(reg_107__in),
    .out(reg_107__out)
  );

  //Wire declarations for instance 'reg_108' (Module coreir_reg)
  wire  reg_108__clk;
  wire [15:0] reg_108__in;
  wire [15:0] reg_108__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_108(
    .clk(reg_108__clk),
    .in(reg_108__in),
    .out(reg_108__out)
  );

  //Wire declarations for instance 'reg_109' (Module coreir_reg)
  wire  reg_109__clk;
  wire [15:0] reg_109__in;
  wire [15:0] reg_109__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_109(
    .clk(reg_109__clk),
    .in(reg_109__in),
    .out(reg_109__out)
  );

  //Wire declarations for instance 'reg_11' (Module coreir_reg)
  wire  reg_11__clk;
  wire [15:0] reg_11__in;
  wire [15:0] reg_11__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_11(
    .clk(reg_11__clk),
    .in(reg_11__in),
    .out(reg_11__out)
  );

  //Wire declarations for instance 'reg_110' (Module coreir_reg)
  wire  reg_110__clk;
  wire [15:0] reg_110__in;
  wire [15:0] reg_110__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_110(
    .clk(reg_110__clk),
    .in(reg_110__in),
    .out(reg_110__out)
  );

  //Wire declarations for instance 'reg_111' (Module coreir_reg)
  wire  reg_111__clk;
  wire [15:0] reg_111__in;
  wire [15:0] reg_111__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_111(
    .clk(reg_111__clk),
    .in(reg_111__in),
    .out(reg_111__out)
  );

  //Wire declarations for instance 'reg_112' (Module coreir_reg)
  wire  reg_112__clk;
  wire [15:0] reg_112__in;
  wire [15:0] reg_112__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_112(
    .clk(reg_112__clk),
    .in(reg_112__in),
    .out(reg_112__out)
  );

  //Wire declarations for instance 'reg_113' (Module coreir_reg)
  wire  reg_113__clk;
  wire [15:0] reg_113__in;
  wire [15:0] reg_113__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_113(
    .clk(reg_113__clk),
    .in(reg_113__in),
    .out(reg_113__out)
  );

  //Wire declarations for instance 'reg_114' (Module coreir_reg)
  wire  reg_114__clk;
  wire [15:0] reg_114__in;
  wire [15:0] reg_114__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_114(
    .clk(reg_114__clk),
    .in(reg_114__in),
    .out(reg_114__out)
  );

  //Wire declarations for instance 'reg_115' (Module coreir_reg)
  wire  reg_115__clk;
  wire [15:0] reg_115__in;
  wire [15:0] reg_115__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_115(
    .clk(reg_115__clk),
    .in(reg_115__in),
    .out(reg_115__out)
  );

  //Wire declarations for instance 'reg_116' (Module coreir_reg)
  wire  reg_116__clk;
  wire [15:0] reg_116__in;
  wire [15:0] reg_116__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_116(
    .clk(reg_116__clk),
    .in(reg_116__in),
    .out(reg_116__out)
  );

  //Wire declarations for instance 'reg_117' (Module coreir_reg)
  wire  reg_117__clk;
  wire [15:0] reg_117__in;
  wire [15:0] reg_117__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_117(
    .clk(reg_117__clk),
    .in(reg_117__in),
    .out(reg_117__out)
  );

  //Wire declarations for instance 'reg_118' (Module coreir_reg)
  wire  reg_118__clk;
  wire [15:0] reg_118__in;
  wire [15:0] reg_118__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_118(
    .clk(reg_118__clk),
    .in(reg_118__in),
    .out(reg_118__out)
  );

  //Wire declarations for instance 'reg_119' (Module coreir_reg)
  wire  reg_119__clk;
  wire [15:0] reg_119__in;
  wire [15:0] reg_119__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_119(
    .clk(reg_119__clk),
    .in(reg_119__in),
    .out(reg_119__out)
  );

  //Wire declarations for instance 'reg_12' (Module coreir_reg)
  wire  reg_12__clk;
  wire [15:0] reg_12__in;
  wire [15:0] reg_12__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_12(
    .clk(reg_12__clk),
    .in(reg_12__in),
    .out(reg_12__out)
  );

  //Wire declarations for instance 'reg_120' (Module coreir_reg)
  wire  reg_120__clk;
  wire [15:0] reg_120__in;
  wire [15:0] reg_120__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_120(
    .clk(reg_120__clk),
    .in(reg_120__in),
    .out(reg_120__out)
  );

  //Wire declarations for instance 'reg_121' (Module coreir_reg)
  wire  reg_121__clk;
  wire [15:0] reg_121__in;
  wire [15:0] reg_121__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_121(
    .clk(reg_121__clk),
    .in(reg_121__in),
    .out(reg_121__out)
  );

  //Wire declarations for instance 'reg_122' (Module coreir_reg)
  wire  reg_122__clk;
  wire [15:0] reg_122__in;
  wire [15:0] reg_122__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_122(
    .clk(reg_122__clk),
    .in(reg_122__in),
    .out(reg_122__out)
  );

  //Wire declarations for instance 'reg_123' (Module coreir_reg)
  wire  reg_123__clk;
  wire [15:0] reg_123__in;
  wire [15:0] reg_123__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_123(
    .clk(reg_123__clk),
    .in(reg_123__in),
    .out(reg_123__out)
  );

  //Wire declarations for instance 'reg_124' (Module coreir_reg)
  wire  reg_124__clk;
  wire [15:0] reg_124__in;
  wire [15:0] reg_124__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_124(
    .clk(reg_124__clk),
    .in(reg_124__in),
    .out(reg_124__out)
  );

  //Wire declarations for instance 'reg_125' (Module coreir_reg)
  wire  reg_125__clk;
  wire [15:0] reg_125__in;
  wire [15:0] reg_125__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_125(
    .clk(reg_125__clk),
    .in(reg_125__in),
    .out(reg_125__out)
  );

  //Wire declarations for instance 'reg_126' (Module coreir_reg)
  wire  reg_126__clk;
  wire [15:0] reg_126__in;
  wire [15:0] reg_126__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_126(
    .clk(reg_126__clk),
    .in(reg_126__in),
    .out(reg_126__out)
  );

  //Wire declarations for instance 'reg_127' (Module coreir_reg)
  wire  reg_127__clk;
  wire [15:0] reg_127__in;
  wire [15:0] reg_127__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_127(
    .clk(reg_127__clk),
    .in(reg_127__in),
    .out(reg_127__out)
  );

  //Wire declarations for instance 'reg_128' (Module coreir_reg)
  wire  reg_128__clk;
  wire [15:0] reg_128__in;
  wire [15:0] reg_128__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_128(
    .clk(reg_128__clk),
    .in(reg_128__in),
    .out(reg_128__out)
  );

  //Wire declarations for instance 'reg_129' (Module coreir_reg)
  wire  reg_129__clk;
  wire [15:0] reg_129__in;
  wire [15:0] reg_129__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_129(
    .clk(reg_129__clk),
    .in(reg_129__in),
    .out(reg_129__out)
  );

  //Wire declarations for instance 'reg_13' (Module coreir_reg)
  wire  reg_13__clk;
  wire [15:0] reg_13__in;
  wire [15:0] reg_13__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_13(
    .clk(reg_13__clk),
    .in(reg_13__in),
    .out(reg_13__out)
  );

  //Wire declarations for instance 'reg_130' (Module coreir_reg)
  wire  reg_130__clk;
  wire [15:0] reg_130__in;
  wire [15:0] reg_130__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_130(
    .clk(reg_130__clk),
    .in(reg_130__in),
    .out(reg_130__out)
  );

  //Wire declarations for instance 'reg_131' (Module coreir_reg)
  wire  reg_131__clk;
  wire [15:0] reg_131__in;
  wire [15:0] reg_131__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_131(
    .clk(reg_131__clk),
    .in(reg_131__in),
    .out(reg_131__out)
  );

  //Wire declarations for instance 'reg_132' (Module coreir_reg)
  wire  reg_132__clk;
  wire [15:0] reg_132__in;
  wire [15:0] reg_132__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_132(
    .clk(reg_132__clk),
    .in(reg_132__in),
    .out(reg_132__out)
  );

  //Wire declarations for instance 'reg_133' (Module coreir_reg)
  wire  reg_133__clk;
  wire [15:0] reg_133__in;
  wire [15:0] reg_133__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_133(
    .clk(reg_133__clk),
    .in(reg_133__in),
    .out(reg_133__out)
  );

  //Wire declarations for instance 'reg_134' (Module coreir_reg)
  wire  reg_134__clk;
  wire [15:0] reg_134__in;
  wire [15:0] reg_134__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_134(
    .clk(reg_134__clk),
    .in(reg_134__in),
    .out(reg_134__out)
  );

  //Wire declarations for instance 'reg_135' (Module coreir_reg)
  wire  reg_135__clk;
  wire [15:0] reg_135__in;
  wire [15:0] reg_135__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_135(
    .clk(reg_135__clk),
    .in(reg_135__in),
    .out(reg_135__out)
  );

  //Wire declarations for instance 'reg_136' (Module coreir_reg)
  wire  reg_136__clk;
  wire [15:0] reg_136__in;
  wire [15:0] reg_136__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_136(
    .clk(reg_136__clk),
    .in(reg_136__in),
    .out(reg_136__out)
  );

  //Wire declarations for instance 'reg_137' (Module coreir_reg)
  wire  reg_137__clk;
  wire [15:0] reg_137__in;
  wire [15:0] reg_137__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_137(
    .clk(reg_137__clk),
    .in(reg_137__in),
    .out(reg_137__out)
  );

  //Wire declarations for instance 'reg_138' (Module coreir_reg)
  wire  reg_138__clk;
  wire [15:0] reg_138__in;
  wire [15:0] reg_138__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_138(
    .clk(reg_138__clk),
    .in(reg_138__in),
    .out(reg_138__out)
  );

  //Wire declarations for instance 'reg_139' (Module coreir_reg)
  wire  reg_139__clk;
  wire [15:0] reg_139__in;
  wire [15:0] reg_139__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_139(
    .clk(reg_139__clk),
    .in(reg_139__in),
    .out(reg_139__out)
  );

  //Wire declarations for instance 'reg_14' (Module coreir_reg)
  wire  reg_14__clk;
  wire [15:0] reg_14__in;
  wire [15:0] reg_14__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_14(
    .clk(reg_14__clk),
    .in(reg_14__in),
    .out(reg_14__out)
  );

  //Wire declarations for instance 'reg_140' (Module coreir_reg)
  wire  reg_140__clk;
  wire [15:0] reg_140__in;
  wire [15:0] reg_140__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_140(
    .clk(reg_140__clk),
    .in(reg_140__in),
    .out(reg_140__out)
  );

  //Wire declarations for instance 'reg_141' (Module coreir_reg)
  wire  reg_141__clk;
  wire [15:0] reg_141__in;
  wire [15:0] reg_141__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_141(
    .clk(reg_141__clk),
    .in(reg_141__in),
    .out(reg_141__out)
  );

  //Wire declarations for instance 'reg_142' (Module coreir_reg)
  wire  reg_142__clk;
  wire [15:0] reg_142__in;
  wire [15:0] reg_142__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_142(
    .clk(reg_142__clk),
    .in(reg_142__in),
    .out(reg_142__out)
  );

  //Wire declarations for instance 'reg_143' (Module coreir_reg)
  wire  reg_143__clk;
  wire [15:0] reg_143__in;
  wire [15:0] reg_143__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_143(
    .clk(reg_143__clk),
    .in(reg_143__in),
    .out(reg_143__out)
  );

  //Wire declarations for instance 'reg_144' (Module coreir_reg)
  wire  reg_144__clk;
  wire [15:0] reg_144__in;
  wire [15:0] reg_144__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_144(
    .clk(reg_144__clk),
    .in(reg_144__in),
    .out(reg_144__out)
  );

  //Wire declarations for instance 'reg_145' (Module coreir_reg)
  wire  reg_145__clk;
  wire [15:0] reg_145__in;
  wire [15:0] reg_145__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_145(
    .clk(reg_145__clk),
    .in(reg_145__in),
    .out(reg_145__out)
  );

  //Wire declarations for instance 'reg_146' (Module coreir_reg)
  wire  reg_146__clk;
  wire [15:0] reg_146__in;
  wire [15:0] reg_146__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_146(
    .clk(reg_146__clk),
    .in(reg_146__in),
    .out(reg_146__out)
  );

  //Wire declarations for instance 'reg_147' (Module coreir_reg)
  wire  reg_147__clk;
  wire [15:0] reg_147__in;
  wire [15:0] reg_147__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_147(
    .clk(reg_147__clk),
    .in(reg_147__in),
    .out(reg_147__out)
  );

  //Wire declarations for instance 'reg_148' (Module coreir_reg)
  wire  reg_148__clk;
  wire [15:0] reg_148__in;
  wire [15:0] reg_148__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_148(
    .clk(reg_148__clk),
    .in(reg_148__in),
    .out(reg_148__out)
  );

  //Wire declarations for instance 'reg_149' (Module coreir_reg)
  wire  reg_149__clk;
  wire [15:0] reg_149__in;
  wire [15:0] reg_149__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_149(
    .clk(reg_149__clk),
    .in(reg_149__in),
    .out(reg_149__out)
  );

  //Wire declarations for instance 'reg_15' (Module coreir_reg)
  wire  reg_15__clk;
  wire [15:0] reg_15__in;
  wire [15:0] reg_15__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_15(
    .clk(reg_15__clk),
    .in(reg_15__in),
    .out(reg_15__out)
  );

  //Wire declarations for instance 'reg_150' (Module coreir_reg)
  wire  reg_150__clk;
  wire [15:0] reg_150__in;
  wire [15:0] reg_150__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_150(
    .clk(reg_150__clk),
    .in(reg_150__in),
    .out(reg_150__out)
  );

  //Wire declarations for instance 'reg_151' (Module coreir_reg)
  wire  reg_151__clk;
  wire [15:0] reg_151__in;
  wire [15:0] reg_151__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_151(
    .clk(reg_151__clk),
    .in(reg_151__in),
    .out(reg_151__out)
  );

  //Wire declarations for instance 'reg_152' (Module coreir_reg)
  wire  reg_152__clk;
  wire [15:0] reg_152__in;
  wire [15:0] reg_152__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_152(
    .clk(reg_152__clk),
    .in(reg_152__in),
    .out(reg_152__out)
  );

  //Wire declarations for instance 'reg_153' (Module coreir_reg)
  wire  reg_153__clk;
  wire [15:0] reg_153__in;
  wire [15:0] reg_153__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_153(
    .clk(reg_153__clk),
    .in(reg_153__in),
    .out(reg_153__out)
  );

  //Wire declarations for instance 'reg_154' (Module coreir_reg)
  wire  reg_154__clk;
  wire [15:0] reg_154__in;
  wire [15:0] reg_154__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_154(
    .clk(reg_154__clk),
    .in(reg_154__in),
    .out(reg_154__out)
  );

  //Wire declarations for instance 'reg_155' (Module coreir_reg)
  wire  reg_155__clk;
  wire [15:0] reg_155__in;
  wire [15:0] reg_155__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_155(
    .clk(reg_155__clk),
    .in(reg_155__in),
    .out(reg_155__out)
  );

  //Wire declarations for instance 'reg_156' (Module coreir_reg)
  wire  reg_156__clk;
  wire [15:0] reg_156__in;
  wire [15:0] reg_156__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_156(
    .clk(reg_156__clk),
    .in(reg_156__in),
    .out(reg_156__out)
  );

  //Wire declarations for instance 'reg_157' (Module coreir_reg)
  wire  reg_157__clk;
  wire [15:0] reg_157__in;
  wire [15:0] reg_157__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_157(
    .clk(reg_157__clk),
    .in(reg_157__in),
    .out(reg_157__out)
  );

  //Wire declarations for instance 'reg_158' (Module coreir_reg)
  wire  reg_158__clk;
  wire [15:0] reg_158__in;
  wire [15:0] reg_158__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_158(
    .clk(reg_158__clk),
    .in(reg_158__in),
    .out(reg_158__out)
  );

  //Wire declarations for instance 'reg_159' (Module coreir_reg)
  wire  reg_159__clk;
  wire [15:0] reg_159__in;
  wire [15:0] reg_159__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_159(
    .clk(reg_159__clk),
    .in(reg_159__in),
    .out(reg_159__out)
  );

  //Wire declarations for instance 'reg_16' (Module coreir_reg)
  wire  reg_16__clk;
  wire [15:0] reg_16__in;
  wire [15:0] reg_16__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_16(
    .clk(reg_16__clk),
    .in(reg_16__in),
    .out(reg_16__out)
  );

  //Wire declarations for instance 'reg_160' (Module coreir_reg)
  wire  reg_160__clk;
  wire [15:0] reg_160__in;
  wire [15:0] reg_160__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_160(
    .clk(reg_160__clk),
    .in(reg_160__in),
    .out(reg_160__out)
  );

  //Wire declarations for instance 'reg_161' (Module coreir_reg)
  wire  reg_161__clk;
  wire [15:0] reg_161__in;
  wire [15:0] reg_161__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_161(
    .clk(reg_161__clk),
    .in(reg_161__in),
    .out(reg_161__out)
  );

  //Wire declarations for instance 'reg_162' (Module coreir_reg)
  wire  reg_162__clk;
  wire [15:0] reg_162__in;
  wire [15:0] reg_162__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_162(
    .clk(reg_162__clk),
    .in(reg_162__in),
    .out(reg_162__out)
  );

  //Wire declarations for instance 'reg_163' (Module coreir_reg)
  wire  reg_163__clk;
  wire [15:0] reg_163__in;
  wire [15:0] reg_163__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_163(
    .clk(reg_163__clk),
    .in(reg_163__in),
    .out(reg_163__out)
  );

  //Wire declarations for instance 'reg_164' (Module coreir_reg)
  wire  reg_164__clk;
  wire [15:0] reg_164__in;
  wire [15:0] reg_164__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_164(
    .clk(reg_164__clk),
    .in(reg_164__in),
    .out(reg_164__out)
  );

  //Wire declarations for instance 'reg_165' (Module coreir_reg)
  wire  reg_165__clk;
  wire [15:0] reg_165__in;
  wire [15:0] reg_165__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_165(
    .clk(reg_165__clk),
    .in(reg_165__in),
    .out(reg_165__out)
  );

  //Wire declarations for instance 'reg_166' (Module coreir_reg)
  wire  reg_166__clk;
  wire [15:0] reg_166__in;
  wire [15:0] reg_166__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_166(
    .clk(reg_166__clk),
    .in(reg_166__in),
    .out(reg_166__out)
  );

  //Wire declarations for instance 'reg_167' (Module coreir_reg)
  wire  reg_167__clk;
  wire [15:0] reg_167__in;
  wire [15:0] reg_167__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_167(
    .clk(reg_167__clk),
    .in(reg_167__in),
    .out(reg_167__out)
  );

  //Wire declarations for instance 'reg_168' (Module coreir_reg)
  wire  reg_168__clk;
  wire [15:0] reg_168__in;
  wire [15:0] reg_168__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_168(
    .clk(reg_168__clk),
    .in(reg_168__in),
    .out(reg_168__out)
  );

  //Wire declarations for instance 'reg_169' (Module coreir_reg)
  wire  reg_169__clk;
  wire [15:0] reg_169__in;
  wire [15:0] reg_169__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_169(
    .clk(reg_169__clk),
    .in(reg_169__in),
    .out(reg_169__out)
  );

  //Wire declarations for instance 'reg_17' (Module coreir_reg)
  wire  reg_17__clk;
  wire [15:0] reg_17__in;
  wire [15:0] reg_17__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_17(
    .clk(reg_17__clk),
    .in(reg_17__in),
    .out(reg_17__out)
  );

  //Wire declarations for instance 'reg_170' (Module coreir_reg)
  wire  reg_170__clk;
  wire [15:0] reg_170__in;
  wire [15:0] reg_170__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_170(
    .clk(reg_170__clk),
    .in(reg_170__in),
    .out(reg_170__out)
  );

  //Wire declarations for instance 'reg_171' (Module coreir_reg)
  wire  reg_171__clk;
  wire [15:0] reg_171__in;
  wire [15:0] reg_171__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_171(
    .clk(reg_171__clk),
    .in(reg_171__in),
    .out(reg_171__out)
  );

  //Wire declarations for instance 'reg_172' (Module coreir_reg)
  wire  reg_172__clk;
  wire [15:0] reg_172__in;
  wire [15:0] reg_172__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_172(
    .clk(reg_172__clk),
    .in(reg_172__in),
    .out(reg_172__out)
  );

  //Wire declarations for instance 'reg_173' (Module coreir_reg)
  wire  reg_173__clk;
  wire [15:0] reg_173__in;
  wire [15:0] reg_173__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_173(
    .clk(reg_173__clk),
    .in(reg_173__in),
    .out(reg_173__out)
  );

  //Wire declarations for instance 'reg_174' (Module coreir_reg)
  wire  reg_174__clk;
  wire [15:0] reg_174__in;
  wire [15:0] reg_174__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_174(
    .clk(reg_174__clk),
    .in(reg_174__in),
    .out(reg_174__out)
  );

  //Wire declarations for instance 'reg_175' (Module coreir_reg)
  wire  reg_175__clk;
  wire [15:0] reg_175__in;
  wire [15:0] reg_175__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_175(
    .clk(reg_175__clk),
    .in(reg_175__in),
    .out(reg_175__out)
  );

  //Wire declarations for instance 'reg_176' (Module coreir_reg)
  wire  reg_176__clk;
  wire [15:0] reg_176__in;
  wire [15:0] reg_176__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_176(
    .clk(reg_176__clk),
    .in(reg_176__in),
    .out(reg_176__out)
  );

  //Wire declarations for instance 'reg_177' (Module coreir_reg)
  wire  reg_177__clk;
  wire [15:0] reg_177__in;
  wire [15:0] reg_177__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_177(
    .clk(reg_177__clk),
    .in(reg_177__in),
    .out(reg_177__out)
  );

  //Wire declarations for instance 'reg_178' (Module coreir_reg)
  wire  reg_178__clk;
  wire [15:0] reg_178__in;
  wire [15:0] reg_178__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_178(
    .clk(reg_178__clk),
    .in(reg_178__in),
    .out(reg_178__out)
  );

  //Wire declarations for instance 'reg_179' (Module coreir_reg)
  wire  reg_179__clk;
  wire [15:0] reg_179__in;
  wire [15:0] reg_179__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_179(
    .clk(reg_179__clk),
    .in(reg_179__in),
    .out(reg_179__out)
  );

  //Wire declarations for instance 'reg_18' (Module coreir_reg)
  wire  reg_18__clk;
  wire [15:0] reg_18__in;
  wire [15:0] reg_18__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_18(
    .clk(reg_18__clk),
    .in(reg_18__in),
    .out(reg_18__out)
  );

  //Wire declarations for instance 'reg_180' (Module coreir_reg)
  wire  reg_180__clk;
  wire [15:0] reg_180__in;
  wire [15:0] reg_180__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_180(
    .clk(reg_180__clk),
    .in(reg_180__in),
    .out(reg_180__out)
  );

  //Wire declarations for instance 'reg_181' (Module coreir_reg)
  wire  reg_181__clk;
  wire [15:0] reg_181__in;
  wire [15:0] reg_181__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_181(
    .clk(reg_181__clk),
    .in(reg_181__in),
    .out(reg_181__out)
  );

  //Wire declarations for instance 'reg_182' (Module coreir_reg)
  wire  reg_182__clk;
  wire [15:0] reg_182__in;
  wire [15:0] reg_182__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_182(
    .clk(reg_182__clk),
    .in(reg_182__in),
    .out(reg_182__out)
  );

  //Wire declarations for instance 'reg_183' (Module coreir_reg)
  wire  reg_183__clk;
  wire [15:0] reg_183__in;
  wire [15:0] reg_183__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_183(
    .clk(reg_183__clk),
    .in(reg_183__in),
    .out(reg_183__out)
  );

  //Wire declarations for instance 'reg_184' (Module coreir_reg)
  wire  reg_184__clk;
  wire [15:0] reg_184__in;
  wire [15:0] reg_184__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_184(
    .clk(reg_184__clk),
    .in(reg_184__in),
    .out(reg_184__out)
  );

  //Wire declarations for instance 'reg_185' (Module coreir_reg)
  wire  reg_185__clk;
  wire [15:0] reg_185__in;
  wire [15:0] reg_185__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_185(
    .clk(reg_185__clk),
    .in(reg_185__in),
    .out(reg_185__out)
  );

  //Wire declarations for instance 'reg_186' (Module coreir_reg)
  wire  reg_186__clk;
  wire [15:0] reg_186__in;
  wire [15:0] reg_186__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_186(
    .clk(reg_186__clk),
    .in(reg_186__in),
    .out(reg_186__out)
  );

  //Wire declarations for instance 'reg_187' (Module coreir_reg)
  wire  reg_187__clk;
  wire [15:0] reg_187__in;
  wire [15:0] reg_187__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_187(
    .clk(reg_187__clk),
    .in(reg_187__in),
    .out(reg_187__out)
  );

  //Wire declarations for instance 'reg_188' (Module coreir_reg)
  wire  reg_188__clk;
  wire [15:0] reg_188__in;
  wire [15:0] reg_188__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_188(
    .clk(reg_188__clk),
    .in(reg_188__in),
    .out(reg_188__out)
  );

  //Wire declarations for instance 'reg_189' (Module coreir_reg)
  wire  reg_189__clk;
  wire [15:0] reg_189__in;
  wire [15:0] reg_189__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_189(
    .clk(reg_189__clk),
    .in(reg_189__in),
    .out(reg_189__out)
  );

  //Wire declarations for instance 'reg_19' (Module coreir_reg)
  wire  reg_19__clk;
  wire [15:0] reg_19__in;
  wire [15:0] reg_19__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_19(
    .clk(reg_19__clk),
    .in(reg_19__in),
    .out(reg_19__out)
  );

  //Wire declarations for instance 'reg_190' (Module coreir_reg)
  wire  reg_190__clk;
  wire [15:0] reg_190__in;
  wire [15:0] reg_190__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_190(
    .clk(reg_190__clk),
    .in(reg_190__in),
    .out(reg_190__out)
  );

  //Wire declarations for instance 'reg_191' (Module coreir_reg)
  wire  reg_191__clk;
  wire [15:0] reg_191__in;
  wire [15:0] reg_191__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_191(
    .clk(reg_191__clk),
    .in(reg_191__in),
    .out(reg_191__out)
  );

  //Wire declarations for instance 'reg_192' (Module coreir_reg)
  wire  reg_192__clk;
  wire [15:0] reg_192__in;
  wire [15:0] reg_192__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_192(
    .clk(reg_192__clk),
    .in(reg_192__in),
    .out(reg_192__out)
  );

  //Wire declarations for instance 'reg_193' (Module coreir_reg)
  wire  reg_193__clk;
  wire [15:0] reg_193__in;
  wire [15:0] reg_193__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_193(
    .clk(reg_193__clk),
    .in(reg_193__in),
    .out(reg_193__out)
  );

  //Wire declarations for instance 'reg_194' (Module coreir_reg)
  wire  reg_194__clk;
  wire [15:0] reg_194__in;
  wire [15:0] reg_194__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_194(
    .clk(reg_194__clk),
    .in(reg_194__in),
    .out(reg_194__out)
  );

  //Wire declarations for instance 'reg_195' (Module coreir_reg)
  wire  reg_195__clk;
  wire [15:0] reg_195__in;
  wire [15:0] reg_195__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_195(
    .clk(reg_195__clk),
    .in(reg_195__in),
    .out(reg_195__out)
  );

  //Wire declarations for instance 'reg_196' (Module coreir_reg)
  wire  reg_196__clk;
  wire [15:0] reg_196__in;
  wire [15:0] reg_196__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_196(
    .clk(reg_196__clk),
    .in(reg_196__in),
    .out(reg_196__out)
  );

  //Wire declarations for instance 'reg_197' (Module coreir_reg)
  wire  reg_197__clk;
  wire [15:0] reg_197__in;
  wire [15:0] reg_197__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_197(
    .clk(reg_197__clk),
    .in(reg_197__in),
    .out(reg_197__out)
  );

  //Wire declarations for instance 'reg_198' (Module coreir_reg)
  wire  reg_198__clk;
  wire [15:0] reg_198__in;
  wire [15:0] reg_198__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_198(
    .clk(reg_198__clk),
    .in(reg_198__in),
    .out(reg_198__out)
  );

  //Wire declarations for instance 'reg_199' (Module coreir_reg)
  wire  reg_199__clk;
  wire [15:0] reg_199__in;
  wire [15:0] reg_199__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_199(
    .clk(reg_199__clk),
    .in(reg_199__in),
    .out(reg_199__out)
  );

  //Wire declarations for instance 'reg_2' (Module coreir_reg)
  wire  reg_2__clk;
  wire [15:0] reg_2__in;
  wire [15:0] reg_2__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_2(
    .clk(reg_2__clk),
    .in(reg_2__in),
    .out(reg_2__out)
  );

  //Wire declarations for instance 'reg_20' (Module coreir_reg)
  wire  reg_20__clk;
  wire [15:0] reg_20__in;
  wire [15:0] reg_20__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_20(
    .clk(reg_20__clk),
    .in(reg_20__in),
    .out(reg_20__out)
  );

  //Wire declarations for instance 'reg_200' (Module coreir_reg)
  wire  reg_200__clk;
  wire [15:0] reg_200__in;
  wire [15:0] reg_200__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_200(
    .clk(reg_200__clk),
    .in(reg_200__in),
    .out(reg_200__out)
  );

  //Wire declarations for instance 'reg_201' (Module coreir_reg)
  wire  reg_201__clk;
  wire [15:0] reg_201__in;
  wire [15:0] reg_201__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_201(
    .clk(reg_201__clk),
    .in(reg_201__in),
    .out(reg_201__out)
  );

  //Wire declarations for instance 'reg_202' (Module coreir_reg)
  wire  reg_202__clk;
  wire [15:0] reg_202__in;
  wire [15:0] reg_202__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_202(
    .clk(reg_202__clk),
    .in(reg_202__in),
    .out(reg_202__out)
  );

  //Wire declarations for instance 'reg_203' (Module coreir_reg)
  wire  reg_203__clk;
  wire [15:0] reg_203__in;
  wire [15:0] reg_203__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_203(
    .clk(reg_203__clk),
    .in(reg_203__in),
    .out(reg_203__out)
  );

  //Wire declarations for instance 'reg_204' (Module coreir_reg)
  wire  reg_204__clk;
  wire [15:0] reg_204__in;
  wire [15:0] reg_204__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_204(
    .clk(reg_204__clk),
    .in(reg_204__in),
    .out(reg_204__out)
  );

  //Wire declarations for instance 'reg_205' (Module coreir_reg)
  wire  reg_205__clk;
  wire [15:0] reg_205__in;
  wire [15:0] reg_205__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_205(
    .clk(reg_205__clk),
    .in(reg_205__in),
    .out(reg_205__out)
  );

  //Wire declarations for instance 'reg_206' (Module coreir_reg)
  wire  reg_206__clk;
  wire [15:0] reg_206__in;
  wire [15:0] reg_206__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_206(
    .clk(reg_206__clk),
    .in(reg_206__in),
    .out(reg_206__out)
  );

  //Wire declarations for instance 'reg_207' (Module coreir_reg)
  wire  reg_207__clk;
  wire [15:0] reg_207__in;
  wire [15:0] reg_207__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_207(
    .clk(reg_207__clk),
    .in(reg_207__in),
    .out(reg_207__out)
  );

  //Wire declarations for instance 'reg_208' (Module coreir_reg)
  wire  reg_208__clk;
  wire [15:0] reg_208__in;
  wire [15:0] reg_208__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_208(
    .clk(reg_208__clk),
    .in(reg_208__in),
    .out(reg_208__out)
  );

  //Wire declarations for instance 'reg_209' (Module coreir_reg)
  wire  reg_209__clk;
  wire [15:0] reg_209__in;
  wire [15:0] reg_209__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_209(
    .clk(reg_209__clk),
    .in(reg_209__in),
    .out(reg_209__out)
  );

  //Wire declarations for instance 'reg_21' (Module coreir_reg)
  wire  reg_21__clk;
  wire [15:0] reg_21__in;
  wire [15:0] reg_21__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_21(
    .clk(reg_21__clk),
    .in(reg_21__in),
    .out(reg_21__out)
  );

  //Wire declarations for instance 'reg_210' (Module coreir_reg)
  wire  reg_210__clk;
  wire [15:0] reg_210__in;
  wire [15:0] reg_210__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_210(
    .clk(reg_210__clk),
    .in(reg_210__in),
    .out(reg_210__out)
  );

  //Wire declarations for instance 'reg_211' (Module coreir_reg)
  wire  reg_211__clk;
  wire [15:0] reg_211__in;
  wire [15:0] reg_211__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_211(
    .clk(reg_211__clk),
    .in(reg_211__in),
    .out(reg_211__out)
  );

  //Wire declarations for instance 'reg_212' (Module coreir_reg)
  wire  reg_212__clk;
  wire [15:0] reg_212__in;
  wire [15:0] reg_212__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_212(
    .clk(reg_212__clk),
    .in(reg_212__in),
    .out(reg_212__out)
  );

  //Wire declarations for instance 'reg_213' (Module coreir_reg)
  wire  reg_213__clk;
  wire [15:0] reg_213__in;
  wire [15:0] reg_213__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_213(
    .clk(reg_213__clk),
    .in(reg_213__in),
    .out(reg_213__out)
  );

  //Wire declarations for instance 'reg_214' (Module coreir_reg)
  wire  reg_214__clk;
  wire [15:0] reg_214__in;
  wire [15:0] reg_214__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_214(
    .clk(reg_214__clk),
    .in(reg_214__in),
    .out(reg_214__out)
  );

  //Wire declarations for instance 'reg_215' (Module coreir_reg)
  wire  reg_215__clk;
  wire [15:0] reg_215__in;
  wire [15:0] reg_215__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_215(
    .clk(reg_215__clk),
    .in(reg_215__in),
    .out(reg_215__out)
  );

  //Wire declarations for instance 'reg_216' (Module coreir_reg)
  wire  reg_216__clk;
  wire [15:0] reg_216__in;
  wire [15:0] reg_216__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_216(
    .clk(reg_216__clk),
    .in(reg_216__in),
    .out(reg_216__out)
  );

  //Wire declarations for instance 'reg_217' (Module coreir_reg)
  wire  reg_217__clk;
  wire [15:0] reg_217__in;
  wire [15:0] reg_217__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_217(
    .clk(reg_217__clk),
    .in(reg_217__in),
    .out(reg_217__out)
  );

  //Wire declarations for instance 'reg_218' (Module coreir_reg)
  wire  reg_218__clk;
  wire [15:0] reg_218__in;
  wire [15:0] reg_218__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_218(
    .clk(reg_218__clk),
    .in(reg_218__in),
    .out(reg_218__out)
  );

  //Wire declarations for instance 'reg_219' (Module coreir_reg)
  wire  reg_219__clk;
  wire [15:0] reg_219__in;
  wire [15:0] reg_219__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_219(
    .clk(reg_219__clk),
    .in(reg_219__in),
    .out(reg_219__out)
  );

  //Wire declarations for instance 'reg_22' (Module coreir_reg)
  wire  reg_22__clk;
  wire [15:0] reg_22__in;
  wire [15:0] reg_22__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_22(
    .clk(reg_22__clk),
    .in(reg_22__in),
    .out(reg_22__out)
  );

  //Wire declarations for instance 'reg_220' (Module coreir_reg)
  wire  reg_220__clk;
  wire [15:0] reg_220__in;
  wire [15:0] reg_220__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_220(
    .clk(reg_220__clk),
    .in(reg_220__in),
    .out(reg_220__out)
  );

  //Wire declarations for instance 'reg_221' (Module coreir_reg)
  wire  reg_221__clk;
  wire [15:0] reg_221__in;
  wire [15:0] reg_221__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_221(
    .clk(reg_221__clk),
    .in(reg_221__in),
    .out(reg_221__out)
  );

  //Wire declarations for instance 'reg_222' (Module coreir_reg)
  wire  reg_222__clk;
  wire [15:0] reg_222__in;
  wire [15:0] reg_222__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_222(
    .clk(reg_222__clk),
    .in(reg_222__in),
    .out(reg_222__out)
  );

  //Wire declarations for instance 'reg_223' (Module coreir_reg)
  wire  reg_223__clk;
  wire [15:0] reg_223__in;
  wire [15:0] reg_223__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_223(
    .clk(reg_223__clk),
    .in(reg_223__in),
    .out(reg_223__out)
  );

  //Wire declarations for instance 'reg_224' (Module coreir_reg)
  wire  reg_224__clk;
  wire [15:0] reg_224__in;
  wire [15:0] reg_224__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_224(
    .clk(reg_224__clk),
    .in(reg_224__in),
    .out(reg_224__out)
  );

  //Wire declarations for instance 'reg_225' (Module coreir_reg)
  wire  reg_225__clk;
  wire [15:0] reg_225__in;
  wire [15:0] reg_225__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_225(
    .clk(reg_225__clk),
    .in(reg_225__in),
    .out(reg_225__out)
  );

  //Wire declarations for instance 'reg_226' (Module coreir_reg)
  wire  reg_226__clk;
  wire [15:0] reg_226__in;
  wire [15:0] reg_226__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_226(
    .clk(reg_226__clk),
    .in(reg_226__in),
    .out(reg_226__out)
  );

  //Wire declarations for instance 'reg_227' (Module coreir_reg)
  wire  reg_227__clk;
  wire [15:0] reg_227__in;
  wire [15:0] reg_227__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_227(
    .clk(reg_227__clk),
    .in(reg_227__in),
    .out(reg_227__out)
  );

  //Wire declarations for instance 'reg_228' (Module coreir_reg)
  wire  reg_228__clk;
  wire [15:0] reg_228__in;
  wire [15:0] reg_228__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_228(
    .clk(reg_228__clk),
    .in(reg_228__in),
    .out(reg_228__out)
  );

  //Wire declarations for instance 'reg_229' (Module coreir_reg)
  wire  reg_229__clk;
  wire [15:0] reg_229__in;
  wire [15:0] reg_229__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_229(
    .clk(reg_229__clk),
    .in(reg_229__in),
    .out(reg_229__out)
  );

  //Wire declarations for instance 'reg_23' (Module coreir_reg)
  wire  reg_23__clk;
  wire [15:0] reg_23__in;
  wire [15:0] reg_23__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_23(
    .clk(reg_23__clk),
    .in(reg_23__in),
    .out(reg_23__out)
  );

  //Wire declarations for instance 'reg_230' (Module coreir_reg)
  wire  reg_230__clk;
  wire [15:0] reg_230__in;
  wire [15:0] reg_230__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_230(
    .clk(reg_230__clk),
    .in(reg_230__in),
    .out(reg_230__out)
  );

  //Wire declarations for instance 'reg_231' (Module coreir_reg)
  wire  reg_231__clk;
  wire [15:0] reg_231__in;
  wire [15:0] reg_231__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_231(
    .clk(reg_231__clk),
    .in(reg_231__in),
    .out(reg_231__out)
  );

  //Wire declarations for instance 'reg_232' (Module coreir_reg)
  wire  reg_232__clk;
  wire [15:0] reg_232__in;
  wire [15:0] reg_232__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_232(
    .clk(reg_232__clk),
    .in(reg_232__in),
    .out(reg_232__out)
  );

  //Wire declarations for instance 'reg_233' (Module coreir_reg)
  wire  reg_233__clk;
  wire [15:0] reg_233__in;
  wire [15:0] reg_233__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_233(
    .clk(reg_233__clk),
    .in(reg_233__in),
    .out(reg_233__out)
  );

  //Wire declarations for instance 'reg_234' (Module coreir_reg)
  wire  reg_234__clk;
  wire [15:0] reg_234__in;
  wire [15:0] reg_234__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_234(
    .clk(reg_234__clk),
    .in(reg_234__in),
    .out(reg_234__out)
  );

  //Wire declarations for instance 'reg_235' (Module coreir_reg)
  wire  reg_235__clk;
  wire [15:0] reg_235__in;
  wire [15:0] reg_235__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_235(
    .clk(reg_235__clk),
    .in(reg_235__in),
    .out(reg_235__out)
  );

  //Wire declarations for instance 'reg_236' (Module coreir_reg)
  wire  reg_236__clk;
  wire [15:0] reg_236__in;
  wire [15:0] reg_236__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_236(
    .clk(reg_236__clk),
    .in(reg_236__in),
    .out(reg_236__out)
  );

  //Wire declarations for instance 'reg_237' (Module coreir_reg)
  wire  reg_237__clk;
  wire [15:0] reg_237__in;
  wire [15:0] reg_237__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_237(
    .clk(reg_237__clk),
    .in(reg_237__in),
    .out(reg_237__out)
  );

  //Wire declarations for instance 'reg_238' (Module coreir_reg)
  wire  reg_238__clk;
  wire [15:0] reg_238__in;
  wire [15:0] reg_238__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_238(
    .clk(reg_238__clk),
    .in(reg_238__in),
    .out(reg_238__out)
  );

  //Wire declarations for instance 'reg_239' (Module coreir_reg)
  wire  reg_239__clk;
  wire [15:0] reg_239__in;
  wire [15:0] reg_239__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_239(
    .clk(reg_239__clk),
    .in(reg_239__in),
    .out(reg_239__out)
  );

  //Wire declarations for instance 'reg_24' (Module coreir_reg)
  wire  reg_24__clk;
  wire [15:0] reg_24__in;
  wire [15:0] reg_24__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_24(
    .clk(reg_24__clk),
    .in(reg_24__in),
    .out(reg_24__out)
  );

  //Wire declarations for instance 'reg_240' (Module coreir_reg)
  wire  reg_240__clk;
  wire [15:0] reg_240__in;
  wire [15:0] reg_240__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_240(
    .clk(reg_240__clk),
    .in(reg_240__in),
    .out(reg_240__out)
  );

  //Wire declarations for instance 'reg_241' (Module coreir_reg)
  wire  reg_241__clk;
  wire [15:0] reg_241__in;
  wire [15:0] reg_241__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_241(
    .clk(reg_241__clk),
    .in(reg_241__in),
    .out(reg_241__out)
  );

  //Wire declarations for instance 'reg_242' (Module coreir_reg)
  wire  reg_242__clk;
  wire [15:0] reg_242__in;
  wire [15:0] reg_242__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_242(
    .clk(reg_242__clk),
    .in(reg_242__in),
    .out(reg_242__out)
  );

  //Wire declarations for instance 'reg_243' (Module coreir_reg)
  wire  reg_243__clk;
  wire [15:0] reg_243__in;
  wire [15:0] reg_243__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_243(
    .clk(reg_243__clk),
    .in(reg_243__in),
    .out(reg_243__out)
  );

  //Wire declarations for instance 'reg_244' (Module coreir_reg)
  wire  reg_244__clk;
  wire [15:0] reg_244__in;
  wire [15:0] reg_244__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_244(
    .clk(reg_244__clk),
    .in(reg_244__in),
    .out(reg_244__out)
  );

  //Wire declarations for instance 'reg_245' (Module coreir_reg)
  wire  reg_245__clk;
  wire [15:0] reg_245__in;
  wire [15:0] reg_245__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_245(
    .clk(reg_245__clk),
    .in(reg_245__in),
    .out(reg_245__out)
  );

  //Wire declarations for instance 'reg_246' (Module coreir_reg)
  wire  reg_246__clk;
  wire [15:0] reg_246__in;
  wire [15:0] reg_246__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_246(
    .clk(reg_246__clk),
    .in(reg_246__in),
    .out(reg_246__out)
  );

  //Wire declarations for instance 'reg_247' (Module coreir_reg)
  wire  reg_247__clk;
  wire [15:0] reg_247__in;
  wire [15:0] reg_247__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_247(
    .clk(reg_247__clk),
    .in(reg_247__in),
    .out(reg_247__out)
  );

  //Wire declarations for instance 'reg_248' (Module coreir_reg)
  wire  reg_248__clk;
  wire [15:0] reg_248__in;
  wire [15:0] reg_248__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_248(
    .clk(reg_248__clk),
    .in(reg_248__in),
    .out(reg_248__out)
  );

  //Wire declarations for instance 'reg_249' (Module coreir_reg)
  wire  reg_249__clk;
  wire [15:0] reg_249__in;
  wire [15:0] reg_249__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_249(
    .clk(reg_249__clk),
    .in(reg_249__in),
    .out(reg_249__out)
  );

  //Wire declarations for instance 'reg_25' (Module coreir_reg)
  wire  reg_25__clk;
  wire [15:0] reg_25__in;
  wire [15:0] reg_25__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_25(
    .clk(reg_25__clk),
    .in(reg_25__in),
    .out(reg_25__out)
  );

  //Wire declarations for instance 'reg_250' (Module coreir_reg)
  wire  reg_250__clk;
  wire [15:0] reg_250__in;
  wire [15:0] reg_250__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_250(
    .clk(reg_250__clk),
    .in(reg_250__in),
    .out(reg_250__out)
  );

  //Wire declarations for instance 'reg_251' (Module coreir_reg)
  wire  reg_251__clk;
  wire [15:0] reg_251__in;
  wire [15:0] reg_251__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_251(
    .clk(reg_251__clk),
    .in(reg_251__in),
    .out(reg_251__out)
  );

  //Wire declarations for instance 'reg_252' (Module coreir_reg)
  wire  reg_252__clk;
  wire [15:0] reg_252__in;
  wire [15:0] reg_252__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_252(
    .clk(reg_252__clk),
    .in(reg_252__in),
    .out(reg_252__out)
  );

  //Wire declarations for instance 'reg_253' (Module coreir_reg)
  wire  reg_253__clk;
  wire [15:0] reg_253__in;
  wire [15:0] reg_253__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_253(
    .clk(reg_253__clk),
    .in(reg_253__in),
    .out(reg_253__out)
  );

  //Wire declarations for instance 'reg_254' (Module coreir_reg)
  wire  reg_254__clk;
  wire [15:0] reg_254__in;
  wire [15:0] reg_254__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_254(
    .clk(reg_254__clk),
    .in(reg_254__in),
    .out(reg_254__out)
  );

  //Wire declarations for instance 'reg_255' (Module coreir_reg)
  wire  reg_255__clk;
  wire [15:0] reg_255__in;
  wire [15:0] reg_255__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_255(
    .clk(reg_255__clk),
    .in(reg_255__in),
    .out(reg_255__out)
  );

  //Wire declarations for instance 'reg_256' (Module coreir_reg)
  wire  reg_256__clk;
  wire [15:0] reg_256__in;
  wire [15:0] reg_256__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_256(
    .clk(reg_256__clk),
    .in(reg_256__in),
    .out(reg_256__out)
  );

  //Wire declarations for instance 'reg_257' (Module coreir_reg)
  wire  reg_257__clk;
  wire [15:0] reg_257__in;
  wire [15:0] reg_257__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_257(
    .clk(reg_257__clk),
    .in(reg_257__in),
    .out(reg_257__out)
  );

  //Wire declarations for instance 'reg_258' (Module coreir_reg)
  wire  reg_258__clk;
  wire [15:0] reg_258__in;
  wire [15:0] reg_258__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_258(
    .clk(reg_258__clk),
    .in(reg_258__in),
    .out(reg_258__out)
  );

  //Wire declarations for instance 'reg_259' (Module coreir_reg)
  wire  reg_259__clk;
  wire [15:0] reg_259__in;
  wire [15:0] reg_259__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_259(
    .clk(reg_259__clk),
    .in(reg_259__in),
    .out(reg_259__out)
  );

  //Wire declarations for instance 'reg_26' (Module coreir_reg)
  wire  reg_26__clk;
  wire [15:0] reg_26__in;
  wire [15:0] reg_26__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_26(
    .clk(reg_26__clk),
    .in(reg_26__in),
    .out(reg_26__out)
  );

  //Wire declarations for instance 'reg_260' (Module coreir_reg)
  wire  reg_260__clk;
  wire [15:0] reg_260__in;
  wire [15:0] reg_260__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_260(
    .clk(reg_260__clk),
    .in(reg_260__in),
    .out(reg_260__out)
  );

  //Wire declarations for instance 'reg_261' (Module coreir_reg)
  wire  reg_261__clk;
  wire [15:0] reg_261__in;
  wire [15:0] reg_261__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_261(
    .clk(reg_261__clk),
    .in(reg_261__in),
    .out(reg_261__out)
  );

  //Wire declarations for instance 'reg_262' (Module coreir_reg)
  wire  reg_262__clk;
  wire [15:0] reg_262__in;
  wire [15:0] reg_262__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_262(
    .clk(reg_262__clk),
    .in(reg_262__in),
    .out(reg_262__out)
  );

  //Wire declarations for instance 'reg_263' (Module coreir_reg)
  wire  reg_263__clk;
  wire [15:0] reg_263__in;
  wire [15:0] reg_263__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_263(
    .clk(reg_263__clk),
    .in(reg_263__in),
    .out(reg_263__out)
  );

  //Wire declarations for instance 'reg_264' (Module coreir_reg)
  wire  reg_264__clk;
  wire [15:0] reg_264__in;
  wire [15:0] reg_264__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_264(
    .clk(reg_264__clk),
    .in(reg_264__in),
    .out(reg_264__out)
  );

  //Wire declarations for instance 'reg_265' (Module coreir_reg)
  wire  reg_265__clk;
  wire [15:0] reg_265__in;
  wire [15:0] reg_265__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_265(
    .clk(reg_265__clk),
    .in(reg_265__in),
    .out(reg_265__out)
  );

  //Wire declarations for instance 'reg_266' (Module coreir_reg)
  wire  reg_266__clk;
  wire [15:0] reg_266__in;
  wire [15:0] reg_266__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_266(
    .clk(reg_266__clk),
    .in(reg_266__in),
    .out(reg_266__out)
  );

  //Wire declarations for instance 'reg_267' (Module coreir_reg)
  wire  reg_267__clk;
  wire [15:0] reg_267__in;
  wire [15:0] reg_267__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_267(
    .clk(reg_267__clk),
    .in(reg_267__in),
    .out(reg_267__out)
  );

  //Wire declarations for instance 'reg_268' (Module coreir_reg)
  wire  reg_268__clk;
  wire [15:0] reg_268__in;
  wire [15:0] reg_268__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_268(
    .clk(reg_268__clk),
    .in(reg_268__in),
    .out(reg_268__out)
  );

  //Wire declarations for instance 'reg_269' (Module coreir_reg)
  wire  reg_269__clk;
  wire [15:0] reg_269__in;
  wire [15:0] reg_269__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_269(
    .clk(reg_269__clk),
    .in(reg_269__in),
    .out(reg_269__out)
  );

  //Wire declarations for instance 'reg_27' (Module coreir_reg)
  wire  reg_27__clk;
  wire [15:0] reg_27__in;
  wire [15:0] reg_27__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_27(
    .clk(reg_27__clk),
    .in(reg_27__in),
    .out(reg_27__out)
  );

  //Wire declarations for instance 'reg_270' (Module coreir_reg)
  wire  reg_270__clk;
  wire [15:0] reg_270__in;
  wire [15:0] reg_270__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_270(
    .clk(reg_270__clk),
    .in(reg_270__in),
    .out(reg_270__out)
  );

  //Wire declarations for instance 'reg_271' (Module coreir_reg)
  wire  reg_271__clk;
  wire [15:0] reg_271__in;
  wire [15:0] reg_271__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_271(
    .clk(reg_271__clk),
    .in(reg_271__in),
    .out(reg_271__out)
  );

  //Wire declarations for instance 'reg_272' (Module coreir_reg)
  wire  reg_272__clk;
  wire [15:0] reg_272__in;
  wire [15:0] reg_272__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_272(
    .clk(reg_272__clk),
    .in(reg_272__in),
    .out(reg_272__out)
  );

  //Wire declarations for instance 'reg_273' (Module coreir_reg)
  wire  reg_273__clk;
  wire [15:0] reg_273__in;
  wire [15:0] reg_273__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_273(
    .clk(reg_273__clk),
    .in(reg_273__in),
    .out(reg_273__out)
  );

  //Wire declarations for instance 'reg_274' (Module coreir_reg)
  wire  reg_274__clk;
  wire [15:0] reg_274__in;
  wire [15:0] reg_274__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_274(
    .clk(reg_274__clk),
    .in(reg_274__in),
    .out(reg_274__out)
  );

  //Wire declarations for instance 'reg_275' (Module coreir_reg)
  wire  reg_275__clk;
  wire [15:0] reg_275__in;
  wire [15:0] reg_275__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_275(
    .clk(reg_275__clk),
    .in(reg_275__in),
    .out(reg_275__out)
  );

  //Wire declarations for instance 'reg_276' (Module coreir_reg)
  wire  reg_276__clk;
  wire [15:0] reg_276__in;
  wire [15:0] reg_276__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_276(
    .clk(reg_276__clk),
    .in(reg_276__in),
    .out(reg_276__out)
  );

  //Wire declarations for instance 'reg_277' (Module coreir_reg)
  wire  reg_277__clk;
  wire [15:0] reg_277__in;
  wire [15:0] reg_277__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_277(
    .clk(reg_277__clk),
    .in(reg_277__in),
    .out(reg_277__out)
  );

  //Wire declarations for instance 'reg_278' (Module coreir_reg)
  wire  reg_278__clk;
  wire [15:0] reg_278__in;
  wire [15:0] reg_278__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_278(
    .clk(reg_278__clk),
    .in(reg_278__in),
    .out(reg_278__out)
  );

  //Wire declarations for instance 'reg_279' (Module coreir_reg)
  wire  reg_279__clk;
  wire [15:0] reg_279__in;
  wire [15:0] reg_279__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_279(
    .clk(reg_279__clk),
    .in(reg_279__in),
    .out(reg_279__out)
  );

  //Wire declarations for instance 'reg_28' (Module coreir_reg)
  wire  reg_28__clk;
  wire [15:0] reg_28__in;
  wire [15:0] reg_28__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_28(
    .clk(reg_28__clk),
    .in(reg_28__in),
    .out(reg_28__out)
  );

  //Wire declarations for instance 'reg_280' (Module coreir_reg)
  wire  reg_280__clk;
  wire [15:0] reg_280__in;
  wire [15:0] reg_280__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_280(
    .clk(reg_280__clk),
    .in(reg_280__in),
    .out(reg_280__out)
  );

  //Wire declarations for instance 'reg_281' (Module coreir_reg)
  wire  reg_281__clk;
  wire [15:0] reg_281__in;
  wire [15:0] reg_281__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_281(
    .clk(reg_281__clk),
    .in(reg_281__in),
    .out(reg_281__out)
  );

  //Wire declarations for instance 'reg_282' (Module coreir_reg)
  wire  reg_282__clk;
  wire [15:0] reg_282__in;
  wire [15:0] reg_282__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_282(
    .clk(reg_282__clk),
    .in(reg_282__in),
    .out(reg_282__out)
  );

  //Wire declarations for instance 'reg_283' (Module coreir_reg)
  wire  reg_283__clk;
  wire [15:0] reg_283__in;
  wire [15:0] reg_283__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_283(
    .clk(reg_283__clk),
    .in(reg_283__in),
    .out(reg_283__out)
  );

  //Wire declarations for instance 'reg_284' (Module coreir_reg)
  wire  reg_284__clk;
  wire [15:0] reg_284__in;
  wire [15:0] reg_284__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_284(
    .clk(reg_284__clk),
    .in(reg_284__in),
    .out(reg_284__out)
  );

  //Wire declarations for instance 'reg_285' (Module coreir_reg)
  wire  reg_285__clk;
  wire [15:0] reg_285__in;
  wire [15:0] reg_285__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_285(
    .clk(reg_285__clk),
    .in(reg_285__in),
    .out(reg_285__out)
  );

  //Wire declarations for instance 'reg_286' (Module coreir_reg)
  wire  reg_286__clk;
  wire [15:0] reg_286__in;
  wire [15:0] reg_286__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_286(
    .clk(reg_286__clk),
    .in(reg_286__in),
    .out(reg_286__out)
  );

  //Wire declarations for instance 'reg_287' (Module coreir_reg)
  wire  reg_287__clk;
  wire [15:0] reg_287__in;
  wire [15:0] reg_287__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_287(
    .clk(reg_287__clk),
    .in(reg_287__in),
    .out(reg_287__out)
  );

  //Wire declarations for instance 'reg_288' (Module coreir_reg)
  wire  reg_288__clk;
  wire [15:0] reg_288__in;
  wire [15:0] reg_288__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_288(
    .clk(reg_288__clk),
    .in(reg_288__in),
    .out(reg_288__out)
  );

  //Wire declarations for instance 'reg_289' (Module coreir_reg)
  wire  reg_289__clk;
  wire [15:0] reg_289__in;
  wire [15:0] reg_289__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_289(
    .clk(reg_289__clk),
    .in(reg_289__in),
    .out(reg_289__out)
  );

  //Wire declarations for instance 'reg_29' (Module coreir_reg)
  wire  reg_29__clk;
  wire [15:0] reg_29__in;
  wire [15:0] reg_29__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_29(
    .clk(reg_29__clk),
    .in(reg_29__in),
    .out(reg_29__out)
  );

  //Wire declarations for instance 'reg_290' (Module coreir_reg)
  wire  reg_290__clk;
  wire [15:0] reg_290__in;
  wire [15:0] reg_290__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_290(
    .clk(reg_290__clk),
    .in(reg_290__in),
    .out(reg_290__out)
  );

  //Wire declarations for instance 'reg_291' (Module coreir_reg)
  wire  reg_291__clk;
  wire [15:0] reg_291__in;
  wire [15:0] reg_291__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_291(
    .clk(reg_291__clk),
    .in(reg_291__in),
    .out(reg_291__out)
  );

  //Wire declarations for instance 'reg_292' (Module coreir_reg)
  wire  reg_292__clk;
  wire [15:0] reg_292__in;
  wire [15:0] reg_292__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_292(
    .clk(reg_292__clk),
    .in(reg_292__in),
    .out(reg_292__out)
  );

  //Wire declarations for instance 'reg_293' (Module coreir_reg)
  wire  reg_293__clk;
  wire [15:0] reg_293__in;
  wire [15:0] reg_293__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_293(
    .clk(reg_293__clk),
    .in(reg_293__in),
    .out(reg_293__out)
  );

  //Wire declarations for instance 'reg_294' (Module coreir_reg)
  wire  reg_294__clk;
  wire [15:0] reg_294__in;
  wire [15:0] reg_294__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_294(
    .clk(reg_294__clk),
    .in(reg_294__in),
    .out(reg_294__out)
  );

  //Wire declarations for instance 'reg_295' (Module coreir_reg)
  wire  reg_295__clk;
  wire [15:0] reg_295__in;
  wire [15:0] reg_295__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_295(
    .clk(reg_295__clk),
    .in(reg_295__in),
    .out(reg_295__out)
  );

  //Wire declarations for instance 'reg_296' (Module coreir_reg)
  wire  reg_296__clk;
  wire [15:0] reg_296__in;
  wire [15:0] reg_296__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_296(
    .clk(reg_296__clk),
    .in(reg_296__in),
    .out(reg_296__out)
  );

  //Wire declarations for instance 'reg_297' (Module coreir_reg)
  wire  reg_297__clk;
  wire [15:0] reg_297__in;
  wire [15:0] reg_297__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_297(
    .clk(reg_297__clk),
    .in(reg_297__in),
    .out(reg_297__out)
  );

  //Wire declarations for instance 'reg_298' (Module coreir_reg)
  wire  reg_298__clk;
  wire [15:0] reg_298__in;
  wire [15:0] reg_298__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_298(
    .clk(reg_298__clk),
    .in(reg_298__in),
    .out(reg_298__out)
  );

  //Wire declarations for instance 'reg_299' (Module coreir_reg)
  wire  reg_299__clk;
  wire [15:0] reg_299__in;
  wire [15:0] reg_299__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_299(
    .clk(reg_299__clk),
    .in(reg_299__in),
    .out(reg_299__out)
  );

  //Wire declarations for instance 'reg_3' (Module coreir_reg)
  wire  reg_3__clk;
  wire [15:0] reg_3__in;
  wire [15:0] reg_3__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_3(
    .clk(reg_3__clk),
    .in(reg_3__in),
    .out(reg_3__out)
  );

  //Wire declarations for instance 'reg_30' (Module coreir_reg)
  wire  reg_30__clk;
  wire [15:0] reg_30__in;
  wire [15:0] reg_30__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_30(
    .clk(reg_30__clk),
    .in(reg_30__in),
    .out(reg_30__out)
  );

  //Wire declarations for instance 'reg_300' (Module coreir_reg)
  wire  reg_300__clk;
  wire [15:0] reg_300__in;
  wire [15:0] reg_300__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_300(
    .clk(reg_300__clk),
    .in(reg_300__in),
    .out(reg_300__out)
  );

  //Wire declarations for instance 'reg_301' (Module coreir_reg)
  wire  reg_301__clk;
  wire [15:0] reg_301__in;
  wire [15:0] reg_301__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_301(
    .clk(reg_301__clk),
    .in(reg_301__in),
    .out(reg_301__out)
  );

  //Wire declarations for instance 'reg_302' (Module coreir_reg)
  wire  reg_302__clk;
  wire [15:0] reg_302__in;
  wire [15:0] reg_302__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_302(
    .clk(reg_302__clk),
    .in(reg_302__in),
    .out(reg_302__out)
  );

  //Wire declarations for instance 'reg_303' (Module coreir_reg)
  wire  reg_303__clk;
  wire [15:0] reg_303__in;
  wire [15:0] reg_303__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_303(
    .clk(reg_303__clk),
    .in(reg_303__in),
    .out(reg_303__out)
  );

  //Wire declarations for instance 'reg_304' (Module coreir_reg)
  wire  reg_304__clk;
  wire [15:0] reg_304__in;
  wire [15:0] reg_304__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_304(
    .clk(reg_304__clk),
    .in(reg_304__in),
    .out(reg_304__out)
  );

  //Wire declarations for instance 'reg_305' (Module coreir_reg)
  wire  reg_305__clk;
  wire [15:0] reg_305__in;
  wire [15:0] reg_305__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_305(
    .clk(reg_305__clk),
    .in(reg_305__in),
    .out(reg_305__out)
  );

  //Wire declarations for instance 'reg_306' (Module coreir_reg)
  wire  reg_306__clk;
  wire [15:0] reg_306__in;
  wire [15:0] reg_306__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_306(
    .clk(reg_306__clk),
    .in(reg_306__in),
    .out(reg_306__out)
  );

  //Wire declarations for instance 'reg_307' (Module coreir_reg)
  wire  reg_307__clk;
  wire [15:0] reg_307__in;
  wire [15:0] reg_307__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_307(
    .clk(reg_307__clk),
    .in(reg_307__in),
    .out(reg_307__out)
  );

  //Wire declarations for instance 'reg_308' (Module coreir_reg)
  wire  reg_308__clk;
  wire [15:0] reg_308__in;
  wire [15:0] reg_308__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_308(
    .clk(reg_308__clk),
    .in(reg_308__in),
    .out(reg_308__out)
  );

  //Wire declarations for instance 'reg_309' (Module coreir_reg)
  wire  reg_309__clk;
  wire [15:0] reg_309__in;
  wire [15:0] reg_309__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_309(
    .clk(reg_309__clk),
    .in(reg_309__in),
    .out(reg_309__out)
  );

  //Wire declarations for instance 'reg_31' (Module coreir_reg)
  wire  reg_31__clk;
  wire [15:0] reg_31__in;
  wire [15:0] reg_31__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_31(
    .clk(reg_31__clk),
    .in(reg_31__in),
    .out(reg_31__out)
  );

  //Wire declarations for instance 'reg_310' (Module coreir_reg)
  wire  reg_310__clk;
  wire [15:0] reg_310__in;
  wire [15:0] reg_310__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_310(
    .clk(reg_310__clk),
    .in(reg_310__in),
    .out(reg_310__out)
  );

  //Wire declarations for instance 'reg_311' (Module coreir_reg)
  wire  reg_311__clk;
  wire [15:0] reg_311__in;
  wire [15:0] reg_311__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_311(
    .clk(reg_311__clk),
    .in(reg_311__in),
    .out(reg_311__out)
  );

  //Wire declarations for instance 'reg_312' (Module coreir_reg)
  wire  reg_312__clk;
  wire [15:0] reg_312__in;
  wire [15:0] reg_312__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_312(
    .clk(reg_312__clk),
    .in(reg_312__in),
    .out(reg_312__out)
  );

  //Wire declarations for instance 'reg_313' (Module coreir_reg)
  wire  reg_313__clk;
  wire [15:0] reg_313__in;
  wire [15:0] reg_313__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_313(
    .clk(reg_313__clk),
    .in(reg_313__in),
    .out(reg_313__out)
  );

  //Wire declarations for instance 'reg_314' (Module coreir_reg)
  wire  reg_314__clk;
  wire [15:0] reg_314__in;
  wire [15:0] reg_314__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_314(
    .clk(reg_314__clk),
    .in(reg_314__in),
    .out(reg_314__out)
  );

  //Wire declarations for instance 'reg_315' (Module coreir_reg)
  wire  reg_315__clk;
  wire [15:0] reg_315__in;
  wire [15:0] reg_315__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_315(
    .clk(reg_315__clk),
    .in(reg_315__in),
    .out(reg_315__out)
  );

  //Wire declarations for instance 'reg_316' (Module coreir_reg)
  wire  reg_316__clk;
  wire [15:0] reg_316__in;
  wire [15:0] reg_316__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_316(
    .clk(reg_316__clk),
    .in(reg_316__in),
    .out(reg_316__out)
  );

  //Wire declarations for instance 'reg_317' (Module coreir_reg)
  wire  reg_317__clk;
  wire [15:0] reg_317__in;
  wire [15:0] reg_317__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_317(
    .clk(reg_317__clk),
    .in(reg_317__in),
    .out(reg_317__out)
  );

  //Wire declarations for instance 'reg_318' (Module coreir_reg)
  wire  reg_318__clk;
  wire [15:0] reg_318__in;
  wire [15:0] reg_318__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_318(
    .clk(reg_318__clk),
    .in(reg_318__in),
    .out(reg_318__out)
  );

  //Wire declarations for instance 'reg_319' (Module coreir_reg)
  wire  reg_319__clk;
  wire [15:0] reg_319__in;
  wire [15:0] reg_319__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_319(
    .clk(reg_319__clk),
    .in(reg_319__in),
    .out(reg_319__out)
  );

  //Wire declarations for instance 'reg_32' (Module coreir_reg)
  wire  reg_32__clk;
  wire [15:0] reg_32__in;
  wire [15:0] reg_32__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_32(
    .clk(reg_32__clk),
    .in(reg_32__in),
    .out(reg_32__out)
  );

  //Wire declarations for instance 'reg_320' (Module coreir_reg)
  wire  reg_320__clk;
  wire [15:0] reg_320__in;
  wire [15:0] reg_320__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_320(
    .clk(reg_320__clk),
    .in(reg_320__in),
    .out(reg_320__out)
  );

  //Wire declarations for instance 'reg_321' (Module coreir_reg)
  wire  reg_321__clk;
  wire [15:0] reg_321__in;
  wire [15:0] reg_321__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_321(
    .clk(reg_321__clk),
    .in(reg_321__in),
    .out(reg_321__out)
  );

  //Wire declarations for instance 'reg_322' (Module coreir_reg)
  wire  reg_322__clk;
  wire [15:0] reg_322__in;
  wire [15:0] reg_322__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_322(
    .clk(reg_322__clk),
    .in(reg_322__in),
    .out(reg_322__out)
  );

  //Wire declarations for instance 'reg_323' (Module coreir_reg)
  wire  reg_323__clk;
  wire [15:0] reg_323__in;
  wire [15:0] reg_323__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_323(
    .clk(reg_323__clk),
    .in(reg_323__in),
    .out(reg_323__out)
  );

  //Wire declarations for instance 'reg_324' (Module coreir_reg)
  wire  reg_324__clk;
  wire [15:0] reg_324__in;
  wire [15:0] reg_324__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_324(
    .clk(reg_324__clk),
    .in(reg_324__in),
    .out(reg_324__out)
  );

  //Wire declarations for instance 'reg_325' (Module coreir_reg)
  wire  reg_325__clk;
  wire [15:0] reg_325__in;
  wire [15:0] reg_325__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_325(
    .clk(reg_325__clk),
    .in(reg_325__in),
    .out(reg_325__out)
  );

  //Wire declarations for instance 'reg_326' (Module coreir_reg)
  wire  reg_326__clk;
  wire [15:0] reg_326__in;
  wire [15:0] reg_326__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_326(
    .clk(reg_326__clk),
    .in(reg_326__in),
    .out(reg_326__out)
  );

  //Wire declarations for instance 'reg_327' (Module coreir_reg)
  wire  reg_327__clk;
  wire [15:0] reg_327__in;
  wire [15:0] reg_327__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_327(
    .clk(reg_327__clk),
    .in(reg_327__in),
    .out(reg_327__out)
  );

  //Wire declarations for instance 'reg_328' (Module coreir_reg)
  wire  reg_328__clk;
  wire [15:0] reg_328__in;
  wire [15:0] reg_328__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_328(
    .clk(reg_328__clk),
    .in(reg_328__in),
    .out(reg_328__out)
  );

  //Wire declarations for instance 'reg_329' (Module coreir_reg)
  wire  reg_329__clk;
  wire [15:0] reg_329__in;
  wire [15:0] reg_329__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_329(
    .clk(reg_329__clk),
    .in(reg_329__in),
    .out(reg_329__out)
  );

  //Wire declarations for instance 'reg_33' (Module coreir_reg)
  wire  reg_33__clk;
  wire [15:0] reg_33__in;
  wire [15:0] reg_33__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_33(
    .clk(reg_33__clk),
    .in(reg_33__in),
    .out(reg_33__out)
  );

  //Wire declarations for instance 'reg_330' (Module coreir_reg)
  wire  reg_330__clk;
  wire [15:0] reg_330__in;
  wire [15:0] reg_330__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_330(
    .clk(reg_330__clk),
    .in(reg_330__in),
    .out(reg_330__out)
  );

  //Wire declarations for instance 'reg_331' (Module coreir_reg)
  wire  reg_331__clk;
  wire [15:0] reg_331__in;
  wire [15:0] reg_331__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_331(
    .clk(reg_331__clk),
    .in(reg_331__in),
    .out(reg_331__out)
  );

  //Wire declarations for instance 'reg_332' (Module coreir_reg)
  wire  reg_332__clk;
  wire [15:0] reg_332__in;
  wire [15:0] reg_332__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_332(
    .clk(reg_332__clk),
    .in(reg_332__in),
    .out(reg_332__out)
  );

  //Wire declarations for instance 'reg_333' (Module coreir_reg)
  wire  reg_333__clk;
  wire [15:0] reg_333__in;
  wire [15:0] reg_333__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_333(
    .clk(reg_333__clk),
    .in(reg_333__in),
    .out(reg_333__out)
  );

  //Wire declarations for instance 'reg_334' (Module coreir_reg)
  wire  reg_334__clk;
  wire [15:0] reg_334__in;
  wire [15:0] reg_334__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_334(
    .clk(reg_334__clk),
    .in(reg_334__in),
    .out(reg_334__out)
  );

  //Wire declarations for instance 'reg_335' (Module coreir_reg)
  wire  reg_335__clk;
  wire [15:0] reg_335__in;
  wire [15:0] reg_335__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_335(
    .clk(reg_335__clk),
    .in(reg_335__in),
    .out(reg_335__out)
  );

  //Wire declarations for instance 'reg_336' (Module coreir_reg)
  wire  reg_336__clk;
  wire [15:0] reg_336__in;
  wire [15:0] reg_336__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_336(
    .clk(reg_336__clk),
    .in(reg_336__in),
    .out(reg_336__out)
  );

  //Wire declarations for instance 'reg_337' (Module coreir_reg)
  wire  reg_337__clk;
  wire [15:0] reg_337__in;
  wire [15:0] reg_337__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_337(
    .clk(reg_337__clk),
    .in(reg_337__in),
    .out(reg_337__out)
  );

  //Wire declarations for instance 'reg_338' (Module coreir_reg)
  wire  reg_338__clk;
  wire [15:0] reg_338__in;
  wire [15:0] reg_338__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_338(
    .clk(reg_338__clk),
    .in(reg_338__in),
    .out(reg_338__out)
  );

  //Wire declarations for instance 'reg_339' (Module coreir_reg)
  wire  reg_339__clk;
  wire [15:0] reg_339__in;
  wire [15:0] reg_339__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_339(
    .clk(reg_339__clk),
    .in(reg_339__in),
    .out(reg_339__out)
  );

  //Wire declarations for instance 'reg_34' (Module coreir_reg)
  wire  reg_34__clk;
  wire [15:0] reg_34__in;
  wire [15:0] reg_34__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_34(
    .clk(reg_34__clk),
    .in(reg_34__in),
    .out(reg_34__out)
  );

  //Wire declarations for instance 'reg_340' (Module coreir_reg)
  wire  reg_340__clk;
  wire [15:0] reg_340__in;
  wire [15:0] reg_340__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_340(
    .clk(reg_340__clk),
    .in(reg_340__in),
    .out(reg_340__out)
  );

  //Wire declarations for instance 'reg_341' (Module coreir_reg)
  wire  reg_341__clk;
  wire [15:0] reg_341__in;
  wire [15:0] reg_341__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_341(
    .clk(reg_341__clk),
    .in(reg_341__in),
    .out(reg_341__out)
  );

  //Wire declarations for instance 'reg_342' (Module coreir_reg)
  wire  reg_342__clk;
  wire [15:0] reg_342__in;
  wire [15:0] reg_342__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_342(
    .clk(reg_342__clk),
    .in(reg_342__in),
    .out(reg_342__out)
  );

  //Wire declarations for instance 'reg_343' (Module coreir_reg)
  wire  reg_343__clk;
  wire [15:0] reg_343__in;
  wire [15:0] reg_343__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_343(
    .clk(reg_343__clk),
    .in(reg_343__in),
    .out(reg_343__out)
  );

  //Wire declarations for instance 'reg_344' (Module coreir_reg)
  wire  reg_344__clk;
  wire [15:0] reg_344__in;
  wire [15:0] reg_344__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_344(
    .clk(reg_344__clk),
    .in(reg_344__in),
    .out(reg_344__out)
  );

  //Wire declarations for instance 'reg_345' (Module coreir_reg)
  wire  reg_345__clk;
  wire [15:0] reg_345__in;
  wire [15:0] reg_345__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_345(
    .clk(reg_345__clk),
    .in(reg_345__in),
    .out(reg_345__out)
  );

  //Wire declarations for instance 'reg_346' (Module coreir_reg)
  wire  reg_346__clk;
  wire [15:0] reg_346__in;
  wire [15:0] reg_346__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_346(
    .clk(reg_346__clk),
    .in(reg_346__in),
    .out(reg_346__out)
  );

  //Wire declarations for instance 'reg_347' (Module coreir_reg)
  wire  reg_347__clk;
  wire [15:0] reg_347__in;
  wire [15:0] reg_347__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_347(
    .clk(reg_347__clk),
    .in(reg_347__in),
    .out(reg_347__out)
  );

  //Wire declarations for instance 'reg_348' (Module coreir_reg)
  wire  reg_348__clk;
  wire [15:0] reg_348__in;
  wire [15:0] reg_348__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_348(
    .clk(reg_348__clk),
    .in(reg_348__in),
    .out(reg_348__out)
  );

  //Wire declarations for instance 'reg_349' (Module coreir_reg)
  wire  reg_349__clk;
  wire [15:0] reg_349__in;
  wire [15:0] reg_349__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_349(
    .clk(reg_349__clk),
    .in(reg_349__in),
    .out(reg_349__out)
  );

  //Wire declarations for instance 'reg_35' (Module coreir_reg)
  wire  reg_35__clk;
  wire [15:0] reg_35__in;
  wire [15:0] reg_35__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_35(
    .clk(reg_35__clk),
    .in(reg_35__in),
    .out(reg_35__out)
  );

  //Wire declarations for instance 'reg_350' (Module coreir_reg)
  wire  reg_350__clk;
  wire [15:0] reg_350__in;
  wire [15:0] reg_350__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_350(
    .clk(reg_350__clk),
    .in(reg_350__in),
    .out(reg_350__out)
  );

  //Wire declarations for instance 'reg_351' (Module coreir_reg)
  wire  reg_351__clk;
  wire [15:0] reg_351__in;
  wire [15:0] reg_351__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_351(
    .clk(reg_351__clk),
    .in(reg_351__in),
    .out(reg_351__out)
  );

  //Wire declarations for instance 'reg_352' (Module coreir_reg)
  wire  reg_352__clk;
  wire [15:0] reg_352__in;
  wire [15:0] reg_352__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_352(
    .clk(reg_352__clk),
    .in(reg_352__in),
    .out(reg_352__out)
  );

  //Wire declarations for instance 'reg_353' (Module coreir_reg)
  wire  reg_353__clk;
  wire [15:0] reg_353__in;
  wire [15:0] reg_353__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_353(
    .clk(reg_353__clk),
    .in(reg_353__in),
    .out(reg_353__out)
  );

  //Wire declarations for instance 'reg_354' (Module coreir_reg)
  wire  reg_354__clk;
  wire [15:0] reg_354__in;
  wire [15:0] reg_354__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_354(
    .clk(reg_354__clk),
    .in(reg_354__in),
    .out(reg_354__out)
  );

  //Wire declarations for instance 'reg_355' (Module coreir_reg)
  wire  reg_355__clk;
  wire [15:0] reg_355__in;
  wire [15:0] reg_355__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_355(
    .clk(reg_355__clk),
    .in(reg_355__in),
    .out(reg_355__out)
  );

  //Wire declarations for instance 'reg_356' (Module coreir_reg)
  wire  reg_356__clk;
  wire [15:0] reg_356__in;
  wire [15:0] reg_356__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_356(
    .clk(reg_356__clk),
    .in(reg_356__in),
    .out(reg_356__out)
  );

  //Wire declarations for instance 'reg_357' (Module coreir_reg)
  wire  reg_357__clk;
  wire [15:0] reg_357__in;
  wire [15:0] reg_357__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_357(
    .clk(reg_357__clk),
    .in(reg_357__in),
    .out(reg_357__out)
  );

  //Wire declarations for instance 'reg_358' (Module coreir_reg)
  wire  reg_358__clk;
  wire [15:0] reg_358__in;
  wire [15:0] reg_358__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_358(
    .clk(reg_358__clk),
    .in(reg_358__in),
    .out(reg_358__out)
  );

  //Wire declarations for instance 'reg_359' (Module coreir_reg)
  wire  reg_359__clk;
  wire [15:0] reg_359__in;
  wire [15:0] reg_359__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_359(
    .clk(reg_359__clk),
    .in(reg_359__in),
    .out(reg_359__out)
  );

  //Wire declarations for instance 'reg_36' (Module coreir_reg)
  wire  reg_36__clk;
  wire [15:0] reg_36__in;
  wire [15:0] reg_36__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_36(
    .clk(reg_36__clk),
    .in(reg_36__in),
    .out(reg_36__out)
  );

  //Wire declarations for instance 'reg_360' (Module coreir_reg)
  wire  reg_360__clk;
  wire [15:0] reg_360__in;
  wire [15:0] reg_360__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_360(
    .clk(reg_360__clk),
    .in(reg_360__in),
    .out(reg_360__out)
  );

  //Wire declarations for instance 'reg_361' (Module coreir_reg)
  wire  reg_361__clk;
  wire [15:0] reg_361__in;
  wire [15:0] reg_361__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_361(
    .clk(reg_361__clk),
    .in(reg_361__in),
    .out(reg_361__out)
  );

  //Wire declarations for instance 'reg_362' (Module coreir_reg)
  wire  reg_362__clk;
  wire [15:0] reg_362__in;
  wire [15:0] reg_362__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_362(
    .clk(reg_362__clk),
    .in(reg_362__in),
    .out(reg_362__out)
  );

  //Wire declarations for instance 'reg_363' (Module coreir_reg)
  wire  reg_363__clk;
  wire [15:0] reg_363__in;
  wire [15:0] reg_363__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_363(
    .clk(reg_363__clk),
    .in(reg_363__in),
    .out(reg_363__out)
  );

  //Wire declarations for instance 'reg_364' (Module coreir_reg)
  wire  reg_364__clk;
  wire [15:0] reg_364__in;
  wire [15:0] reg_364__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_364(
    .clk(reg_364__clk),
    .in(reg_364__in),
    .out(reg_364__out)
  );

  //Wire declarations for instance 'reg_365' (Module coreir_reg)
  wire  reg_365__clk;
  wire [15:0] reg_365__in;
  wire [15:0] reg_365__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_365(
    .clk(reg_365__clk),
    .in(reg_365__in),
    .out(reg_365__out)
  );

  //Wire declarations for instance 'reg_366' (Module coreir_reg)
  wire  reg_366__clk;
  wire [15:0] reg_366__in;
  wire [15:0] reg_366__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_366(
    .clk(reg_366__clk),
    .in(reg_366__in),
    .out(reg_366__out)
  );

  //Wire declarations for instance 'reg_367' (Module coreir_reg)
  wire  reg_367__clk;
  wire [15:0] reg_367__in;
  wire [15:0] reg_367__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_367(
    .clk(reg_367__clk),
    .in(reg_367__in),
    .out(reg_367__out)
  );

  //Wire declarations for instance 'reg_368' (Module coreir_reg)
  wire  reg_368__clk;
  wire [15:0] reg_368__in;
  wire [15:0] reg_368__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_368(
    .clk(reg_368__clk),
    .in(reg_368__in),
    .out(reg_368__out)
  );

  //Wire declarations for instance 'reg_369' (Module coreir_reg)
  wire  reg_369__clk;
  wire [15:0] reg_369__in;
  wire [15:0] reg_369__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_369(
    .clk(reg_369__clk),
    .in(reg_369__in),
    .out(reg_369__out)
  );

  //Wire declarations for instance 'reg_37' (Module coreir_reg)
  wire  reg_37__clk;
  wire [15:0] reg_37__in;
  wire [15:0] reg_37__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_37(
    .clk(reg_37__clk),
    .in(reg_37__in),
    .out(reg_37__out)
  );

  //Wire declarations for instance 'reg_370' (Module coreir_reg)
  wire  reg_370__clk;
  wire [15:0] reg_370__in;
  wire [15:0] reg_370__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_370(
    .clk(reg_370__clk),
    .in(reg_370__in),
    .out(reg_370__out)
  );

  //Wire declarations for instance 'reg_371' (Module coreir_reg)
  wire  reg_371__clk;
  wire [15:0] reg_371__in;
  wire [15:0] reg_371__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_371(
    .clk(reg_371__clk),
    .in(reg_371__in),
    .out(reg_371__out)
  );

  //Wire declarations for instance 'reg_372' (Module coreir_reg)
  wire  reg_372__clk;
  wire [15:0] reg_372__in;
  wire [15:0] reg_372__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_372(
    .clk(reg_372__clk),
    .in(reg_372__in),
    .out(reg_372__out)
  );

  //Wire declarations for instance 'reg_373' (Module coreir_reg)
  wire  reg_373__clk;
  wire [15:0] reg_373__in;
  wire [15:0] reg_373__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_373(
    .clk(reg_373__clk),
    .in(reg_373__in),
    .out(reg_373__out)
  );

  //Wire declarations for instance 'reg_374' (Module coreir_reg)
  wire  reg_374__clk;
  wire [15:0] reg_374__in;
  wire [15:0] reg_374__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_374(
    .clk(reg_374__clk),
    .in(reg_374__in),
    .out(reg_374__out)
  );

  //Wire declarations for instance 'reg_375' (Module coreir_reg)
  wire  reg_375__clk;
  wire [15:0] reg_375__in;
  wire [15:0] reg_375__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_375(
    .clk(reg_375__clk),
    .in(reg_375__in),
    .out(reg_375__out)
  );

  //Wire declarations for instance 'reg_376' (Module coreir_reg)
  wire  reg_376__clk;
  wire [15:0] reg_376__in;
  wire [15:0] reg_376__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_376(
    .clk(reg_376__clk),
    .in(reg_376__in),
    .out(reg_376__out)
  );

  //Wire declarations for instance 'reg_377' (Module coreir_reg)
  wire  reg_377__clk;
  wire [15:0] reg_377__in;
  wire [15:0] reg_377__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_377(
    .clk(reg_377__clk),
    .in(reg_377__in),
    .out(reg_377__out)
  );

  //Wire declarations for instance 'reg_378' (Module coreir_reg)
  wire  reg_378__clk;
  wire [15:0] reg_378__in;
  wire [15:0] reg_378__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_378(
    .clk(reg_378__clk),
    .in(reg_378__in),
    .out(reg_378__out)
  );

  //Wire declarations for instance 'reg_379' (Module coreir_reg)
  wire  reg_379__clk;
  wire [15:0] reg_379__in;
  wire [15:0] reg_379__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_379(
    .clk(reg_379__clk),
    .in(reg_379__in),
    .out(reg_379__out)
  );

  //Wire declarations for instance 'reg_38' (Module coreir_reg)
  wire  reg_38__clk;
  wire [15:0] reg_38__in;
  wire [15:0] reg_38__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_38(
    .clk(reg_38__clk),
    .in(reg_38__in),
    .out(reg_38__out)
  );

  //Wire declarations for instance 'reg_380' (Module coreir_reg)
  wire  reg_380__clk;
  wire [15:0] reg_380__in;
  wire [15:0] reg_380__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_380(
    .clk(reg_380__clk),
    .in(reg_380__in),
    .out(reg_380__out)
  );

  //Wire declarations for instance 'reg_381' (Module coreir_reg)
  wire  reg_381__clk;
  wire [15:0] reg_381__in;
  wire [15:0] reg_381__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_381(
    .clk(reg_381__clk),
    .in(reg_381__in),
    .out(reg_381__out)
  );

  //Wire declarations for instance 'reg_382' (Module coreir_reg)
  wire  reg_382__clk;
  wire [15:0] reg_382__in;
  wire [15:0] reg_382__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_382(
    .clk(reg_382__clk),
    .in(reg_382__in),
    .out(reg_382__out)
  );

  //Wire declarations for instance 'reg_383' (Module coreir_reg)
  wire  reg_383__clk;
  wire [15:0] reg_383__in;
  wire [15:0] reg_383__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_383(
    .clk(reg_383__clk),
    .in(reg_383__in),
    .out(reg_383__out)
  );

  //Wire declarations for instance 'reg_384' (Module coreir_reg)
  wire  reg_384__clk;
  wire [15:0] reg_384__in;
  wire [15:0] reg_384__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_384(
    .clk(reg_384__clk),
    .in(reg_384__in),
    .out(reg_384__out)
  );

  //Wire declarations for instance 'reg_385' (Module coreir_reg)
  wire  reg_385__clk;
  wire [15:0] reg_385__in;
  wire [15:0] reg_385__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_385(
    .clk(reg_385__clk),
    .in(reg_385__in),
    .out(reg_385__out)
  );

  //Wire declarations for instance 'reg_386' (Module coreir_reg)
  wire  reg_386__clk;
  wire [15:0] reg_386__in;
  wire [15:0] reg_386__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_386(
    .clk(reg_386__clk),
    .in(reg_386__in),
    .out(reg_386__out)
  );

  //Wire declarations for instance 'reg_387' (Module coreir_reg)
  wire  reg_387__clk;
  wire [15:0] reg_387__in;
  wire [15:0] reg_387__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_387(
    .clk(reg_387__clk),
    .in(reg_387__in),
    .out(reg_387__out)
  );

  //Wire declarations for instance 'reg_388' (Module coreir_reg)
  wire  reg_388__clk;
  wire [15:0] reg_388__in;
  wire [15:0] reg_388__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_388(
    .clk(reg_388__clk),
    .in(reg_388__in),
    .out(reg_388__out)
  );

  //Wire declarations for instance 'reg_389' (Module coreir_reg)
  wire  reg_389__clk;
  wire [15:0] reg_389__in;
  wire [15:0] reg_389__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_389(
    .clk(reg_389__clk),
    .in(reg_389__in),
    .out(reg_389__out)
  );

  //Wire declarations for instance 'reg_39' (Module coreir_reg)
  wire  reg_39__clk;
  wire [15:0] reg_39__in;
  wire [15:0] reg_39__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_39(
    .clk(reg_39__clk),
    .in(reg_39__in),
    .out(reg_39__out)
  );

  //Wire declarations for instance 'reg_390' (Module coreir_reg)
  wire  reg_390__clk;
  wire [15:0] reg_390__in;
  wire [15:0] reg_390__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_390(
    .clk(reg_390__clk),
    .in(reg_390__in),
    .out(reg_390__out)
  );

  //Wire declarations for instance 'reg_391' (Module coreir_reg)
  wire  reg_391__clk;
  wire [15:0] reg_391__in;
  wire [15:0] reg_391__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_391(
    .clk(reg_391__clk),
    .in(reg_391__in),
    .out(reg_391__out)
  );

  //Wire declarations for instance 'reg_392' (Module coreir_reg)
  wire  reg_392__clk;
  wire [15:0] reg_392__in;
  wire [15:0] reg_392__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_392(
    .clk(reg_392__clk),
    .in(reg_392__in),
    .out(reg_392__out)
  );

  //Wire declarations for instance 'reg_393' (Module coreir_reg)
  wire  reg_393__clk;
  wire [15:0] reg_393__in;
  wire [15:0] reg_393__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_393(
    .clk(reg_393__clk),
    .in(reg_393__in),
    .out(reg_393__out)
  );

  //Wire declarations for instance 'reg_394' (Module coreir_reg)
  wire  reg_394__clk;
  wire [15:0] reg_394__in;
  wire [15:0] reg_394__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_394(
    .clk(reg_394__clk),
    .in(reg_394__in),
    .out(reg_394__out)
  );

  //Wire declarations for instance 'reg_395' (Module coreir_reg)
  wire  reg_395__clk;
  wire [15:0] reg_395__in;
  wire [15:0] reg_395__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_395(
    .clk(reg_395__clk),
    .in(reg_395__in),
    .out(reg_395__out)
  );

  //Wire declarations for instance 'reg_396' (Module coreir_reg)
  wire  reg_396__clk;
  wire [15:0] reg_396__in;
  wire [15:0] reg_396__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_396(
    .clk(reg_396__clk),
    .in(reg_396__in),
    .out(reg_396__out)
  );

  //Wire declarations for instance 'reg_397' (Module coreir_reg)
  wire  reg_397__clk;
  wire [15:0] reg_397__in;
  wire [15:0] reg_397__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_397(
    .clk(reg_397__clk),
    .in(reg_397__in),
    .out(reg_397__out)
  );

  //Wire declarations for instance 'reg_398' (Module coreir_reg)
  wire  reg_398__clk;
  wire [15:0] reg_398__in;
  wire [15:0] reg_398__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_398(
    .clk(reg_398__clk),
    .in(reg_398__in),
    .out(reg_398__out)
  );

  //Wire declarations for instance 'reg_399' (Module coreir_reg)
  wire  reg_399__clk;
  wire [15:0] reg_399__in;
  wire [15:0] reg_399__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_399(
    .clk(reg_399__clk),
    .in(reg_399__in),
    .out(reg_399__out)
  );

  //Wire declarations for instance 'reg_4' (Module coreir_reg)
  wire  reg_4__clk;
  wire [15:0] reg_4__in;
  wire [15:0] reg_4__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_4(
    .clk(reg_4__clk),
    .in(reg_4__in),
    .out(reg_4__out)
  );

  //Wire declarations for instance 'reg_40' (Module coreir_reg)
  wire  reg_40__clk;
  wire [15:0] reg_40__in;
  wire [15:0] reg_40__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_40(
    .clk(reg_40__clk),
    .in(reg_40__in),
    .out(reg_40__out)
  );

  //Wire declarations for instance 'reg_400' (Module coreir_reg)
  wire  reg_400__clk;
  wire [15:0] reg_400__in;
  wire [15:0] reg_400__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_400(
    .clk(reg_400__clk),
    .in(reg_400__in),
    .out(reg_400__out)
  );

  //Wire declarations for instance 'reg_401' (Module coreir_reg)
  wire  reg_401__clk;
  wire [15:0] reg_401__in;
  wire [15:0] reg_401__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_401(
    .clk(reg_401__clk),
    .in(reg_401__in),
    .out(reg_401__out)
  );

  //Wire declarations for instance 'reg_402' (Module coreir_reg)
  wire  reg_402__clk;
  wire [15:0] reg_402__in;
  wire [15:0] reg_402__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_402(
    .clk(reg_402__clk),
    .in(reg_402__in),
    .out(reg_402__out)
  );

  //Wire declarations for instance 'reg_403' (Module coreir_reg)
  wire  reg_403__clk;
  wire [15:0] reg_403__in;
  wire [15:0] reg_403__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_403(
    .clk(reg_403__clk),
    .in(reg_403__in),
    .out(reg_403__out)
  );

  //Wire declarations for instance 'reg_404' (Module coreir_reg)
  wire  reg_404__clk;
  wire [15:0] reg_404__in;
  wire [15:0] reg_404__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_404(
    .clk(reg_404__clk),
    .in(reg_404__in),
    .out(reg_404__out)
  );

  //Wire declarations for instance 'reg_405' (Module coreir_reg)
  wire  reg_405__clk;
  wire [15:0] reg_405__in;
  wire [15:0] reg_405__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_405(
    .clk(reg_405__clk),
    .in(reg_405__in),
    .out(reg_405__out)
  );

  //Wire declarations for instance 'reg_406' (Module coreir_reg)
  wire  reg_406__clk;
  wire [15:0] reg_406__in;
  wire [15:0] reg_406__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_406(
    .clk(reg_406__clk),
    .in(reg_406__in),
    .out(reg_406__out)
  );

  //Wire declarations for instance 'reg_407' (Module coreir_reg)
  wire  reg_407__clk;
  wire [15:0] reg_407__in;
  wire [15:0] reg_407__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_407(
    .clk(reg_407__clk),
    .in(reg_407__in),
    .out(reg_407__out)
  );

  //Wire declarations for instance 'reg_408' (Module coreir_reg)
  wire  reg_408__clk;
  wire [15:0] reg_408__in;
  wire [15:0] reg_408__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_408(
    .clk(reg_408__clk),
    .in(reg_408__in),
    .out(reg_408__out)
  );

  //Wire declarations for instance 'reg_409' (Module coreir_reg)
  wire  reg_409__clk;
  wire [15:0] reg_409__in;
  wire [15:0] reg_409__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_409(
    .clk(reg_409__clk),
    .in(reg_409__in),
    .out(reg_409__out)
  );

  //Wire declarations for instance 'reg_41' (Module coreir_reg)
  wire  reg_41__clk;
  wire [15:0] reg_41__in;
  wire [15:0] reg_41__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_41(
    .clk(reg_41__clk),
    .in(reg_41__in),
    .out(reg_41__out)
  );

  //Wire declarations for instance 'reg_410' (Module coreir_reg)
  wire  reg_410__clk;
  wire [15:0] reg_410__in;
  wire [15:0] reg_410__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_410(
    .clk(reg_410__clk),
    .in(reg_410__in),
    .out(reg_410__out)
  );

  //Wire declarations for instance 'reg_411' (Module coreir_reg)
  wire  reg_411__clk;
  wire [15:0] reg_411__in;
  wire [15:0] reg_411__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_411(
    .clk(reg_411__clk),
    .in(reg_411__in),
    .out(reg_411__out)
  );

  //Wire declarations for instance 'reg_412' (Module coreir_reg)
  wire  reg_412__clk;
  wire [15:0] reg_412__in;
  wire [15:0] reg_412__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_412(
    .clk(reg_412__clk),
    .in(reg_412__in),
    .out(reg_412__out)
  );

  //Wire declarations for instance 'reg_413' (Module coreir_reg)
  wire  reg_413__clk;
  wire [15:0] reg_413__in;
  wire [15:0] reg_413__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_413(
    .clk(reg_413__clk),
    .in(reg_413__in),
    .out(reg_413__out)
  );

  //Wire declarations for instance 'reg_414' (Module coreir_reg)
  wire  reg_414__clk;
  wire [15:0] reg_414__in;
  wire [15:0] reg_414__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_414(
    .clk(reg_414__clk),
    .in(reg_414__in),
    .out(reg_414__out)
  );

  //Wire declarations for instance 'reg_415' (Module coreir_reg)
  wire  reg_415__clk;
  wire [15:0] reg_415__in;
  wire [15:0] reg_415__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_415(
    .clk(reg_415__clk),
    .in(reg_415__in),
    .out(reg_415__out)
  );

  //Wire declarations for instance 'reg_416' (Module coreir_reg)
  wire  reg_416__clk;
  wire [15:0] reg_416__in;
  wire [15:0] reg_416__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_416(
    .clk(reg_416__clk),
    .in(reg_416__in),
    .out(reg_416__out)
  );

  //Wire declarations for instance 'reg_417' (Module coreir_reg)
  wire  reg_417__clk;
  wire [15:0] reg_417__in;
  wire [15:0] reg_417__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_417(
    .clk(reg_417__clk),
    .in(reg_417__in),
    .out(reg_417__out)
  );

  //Wire declarations for instance 'reg_418' (Module coreir_reg)
  wire  reg_418__clk;
  wire [15:0] reg_418__in;
  wire [15:0] reg_418__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_418(
    .clk(reg_418__clk),
    .in(reg_418__in),
    .out(reg_418__out)
  );

  //Wire declarations for instance 'reg_419' (Module coreir_reg)
  wire  reg_419__clk;
  wire [15:0] reg_419__in;
  wire [15:0] reg_419__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_419(
    .clk(reg_419__clk),
    .in(reg_419__in),
    .out(reg_419__out)
  );

  //Wire declarations for instance 'reg_42' (Module coreir_reg)
  wire  reg_42__clk;
  wire [15:0] reg_42__in;
  wire [15:0] reg_42__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_42(
    .clk(reg_42__clk),
    .in(reg_42__in),
    .out(reg_42__out)
  );

  //Wire declarations for instance 'reg_420' (Module coreir_reg)
  wire  reg_420__clk;
  wire [15:0] reg_420__in;
  wire [15:0] reg_420__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_420(
    .clk(reg_420__clk),
    .in(reg_420__in),
    .out(reg_420__out)
  );

  //Wire declarations for instance 'reg_421' (Module coreir_reg)
  wire  reg_421__clk;
  wire [15:0] reg_421__in;
  wire [15:0] reg_421__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_421(
    .clk(reg_421__clk),
    .in(reg_421__in),
    .out(reg_421__out)
  );

  //Wire declarations for instance 'reg_422' (Module coreir_reg)
  wire  reg_422__clk;
  wire [15:0] reg_422__in;
  wire [15:0] reg_422__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_422(
    .clk(reg_422__clk),
    .in(reg_422__in),
    .out(reg_422__out)
  );

  //Wire declarations for instance 'reg_423' (Module coreir_reg)
  wire  reg_423__clk;
  wire [15:0] reg_423__in;
  wire [15:0] reg_423__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_423(
    .clk(reg_423__clk),
    .in(reg_423__in),
    .out(reg_423__out)
  );

  //Wire declarations for instance 'reg_424' (Module coreir_reg)
  wire  reg_424__clk;
  wire [15:0] reg_424__in;
  wire [15:0] reg_424__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_424(
    .clk(reg_424__clk),
    .in(reg_424__in),
    .out(reg_424__out)
  );

  //Wire declarations for instance 'reg_425' (Module coreir_reg)
  wire  reg_425__clk;
  wire [15:0] reg_425__in;
  wire [15:0] reg_425__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_425(
    .clk(reg_425__clk),
    .in(reg_425__in),
    .out(reg_425__out)
  );

  //Wire declarations for instance 'reg_426' (Module coreir_reg)
  wire  reg_426__clk;
  wire [15:0] reg_426__in;
  wire [15:0] reg_426__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_426(
    .clk(reg_426__clk),
    .in(reg_426__in),
    .out(reg_426__out)
  );

  //Wire declarations for instance 'reg_427' (Module coreir_reg)
  wire  reg_427__clk;
  wire [15:0] reg_427__in;
  wire [15:0] reg_427__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_427(
    .clk(reg_427__clk),
    .in(reg_427__in),
    .out(reg_427__out)
  );

  //Wire declarations for instance 'reg_428' (Module coreir_reg)
  wire  reg_428__clk;
  wire [15:0] reg_428__in;
  wire [15:0] reg_428__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_428(
    .clk(reg_428__clk),
    .in(reg_428__in),
    .out(reg_428__out)
  );

  //Wire declarations for instance 'reg_429' (Module coreir_reg)
  wire  reg_429__clk;
  wire [15:0] reg_429__in;
  wire [15:0] reg_429__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_429(
    .clk(reg_429__clk),
    .in(reg_429__in),
    .out(reg_429__out)
  );

  //Wire declarations for instance 'reg_43' (Module coreir_reg)
  wire  reg_43__clk;
  wire [15:0] reg_43__in;
  wire [15:0] reg_43__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_43(
    .clk(reg_43__clk),
    .in(reg_43__in),
    .out(reg_43__out)
  );

  //Wire declarations for instance 'reg_430' (Module coreir_reg)
  wire  reg_430__clk;
  wire [15:0] reg_430__in;
  wire [15:0] reg_430__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_430(
    .clk(reg_430__clk),
    .in(reg_430__in),
    .out(reg_430__out)
  );

  //Wire declarations for instance 'reg_431' (Module coreir_reg)
  wire  reg_431__clk;
  wire [15:0] reg_431__in;
  wire [15:0] reg_431__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_431(
    .clk(reg_431__clk),
    .in(reg_431__in),
    .out(reg_431__out)
  );

  //Wire declarations for instance 'reg_432' (Module coreir_reg)
  wire  reg_432__clk;
  wire [15:0] reg_432__in;
  wire [15:0] reg_432__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_432(
    .clk(reg_432__clk),
    .in(reg_432__in),
    .out(reg_432__out)
  );

  //Wire declarations for instance 'reg_433' (Module coreir_reg)
  wire  reg_433__clk;
  wire [15:0] reg_433__in;
  wire [15:0] reg_433__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_433(
    .clk(reg_433__clk),
    .in(reg_433__in),
    .out(reg_433__out)
  );

  //Wire declarations for instance 'reg_434' (Module coreir_reg)
  wire  reg_434__clk;
  wire [15:0] reg_434__in;
  wire [15:0] reg_434__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_434(
    .clk(reg_434__clk),
    .in(reg_434__in),
    .out(reg_434__out)
  );

  //Wire declarations for instance 'reg_435' (Module coreir_reg)
  wire  reg_435__clk;
  wire [15:0] reg_435__in;
  wire [15:0] reg_435__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_435(
    .clk(reg_435__clk),
    .in(reg_435__in),
    .out(reg_435__out)
  );

  //Wire declarations for instance 'reg_436' (Module coreir_reg)
  wire  reg_436__clk;
  wire [15:0] reg_436__in;
  wire [15:0] reg_436__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_436(
    .clk(reg_436__clk),
    .in(reg_436__in),
    .out(reg_436__out)
  );

  //Wire declarations for instance 'reg_437' (Module coreir_reg)
  wire  reg_437__clk;
  wire [15:0] reg_437__in;
  wire [15:0] reg_437__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_437(
    .clk(reg_437__clk),
    .in(reg_437__in),
    .out(reg_437__out)
  );

  //Wire declarations for instance 'reg_438' (Module coreir_reg)
  wire  reg_438__clk;
  wire [15:0] reg_438__in;
  wire [15:0] reg_438__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_438(
    .clk(reg_438__clk),
    .in(reg_438__in),
    .out(reg_438__out)
  );

  //Wire declarations for instance 'reg_439' (Module coreir_reg)
  wire  reg_439__clk;
  wire [15:0] reg_439__in;
  wire [15:0] reg_439__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_439(
    .clk(reg_439__clk),
    .in(reg_439__in),
    .out(reg_439__out)
  );

  //Wire declarations for instance 'reg_44' (Module coreir_reg)
  wire  reg_44__clk;
  wire [15:0] reg_44__in;
  wire [15:0] reg_44__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_44(
    .clk(reg_44__clk),
    .in(reg_44__in),
    .out(reg_44__out)
  );

  //Wire declarations for instance 'reg_440' (Module coreir_reg)
  wire  reg_440__clk;
  wire [15:0] reg_440__in;
  wire [15:0] reg_440__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_440(
    .clk(reg_440__clk),
    .in(reg_440__in),
    .out(reg_440__out)
  );

  //Wire declarations for instance 'reg_441' (Module coreir_reg)
  wire  reg_441__clk;
  wire [15:0] reg_441__in;
  wire [15:0] reg_441__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_441(
    .clk(reg_441__clk),
    .in(reg_441__in),
    .out(reg_441__out)
  );

  //Wire declarations for instance 'reg_442' (Module coreir_reg)
  wire  reg_442__clk;
  wire [15:0] reg_442__in;
  wire [15:0] reg_442__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_442(
    .clk(reg_442__clk),
    .in(reg_442__in),
    .out(reg_442__out)
  );

  //Wire declarations for instance 'reg_443' (Module coreir_reg)
  wire  reg_443__clk;
  wire [15:0] reg_443__in;
  wire [15:0] reg_443__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_443(
    .clk(reg_443__clk),
    .in(reg_443__in),
    .out(reg_443__out)
  );

  //Wire declarations for instance 'reg_444' (Module coreir_reg)
  wire  reg_444__clk;
  wire [15:0] reg_444__in;
  wire [15:0] reg_444__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_444(
    .clk(reg_444__clk),
    .in(reg_444__in),
    .out(reg_444__out)
  );

  //Wire declarations for instance 'reg_445' (Module coreir_reg)
  wire  reg_445__clk;
  wire [15:0] reg_445__in;
  wire [15:0] reg_445__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_445(
    .clk(reg_445__clk),
    .in(reg_445__in),
    .out(reg_445__out)
  );

  //Wire declarations for instance 'reg_446' (Module coreir_reg)
  wire  reg_446__clk;
  wire [15:0] reg_446__in;
  wire [15:0] reg_446__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_446(
    .clk(reg_446__clk),
    .in(reg_446__in),
    .out(reg_446__out)
  );

  //Wire declarations for instance 'reg_447' (Module coreir_reg)
  wire  reg_447__clk;
  wire [15:0] reg_447__in;
  wire [15:0] reg_447__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_447(
    .clk(reg_447__clk),
    .in(reg_447__in),
    .out(reg_447__out)
  );

  //Wire declarations for instance 'reg_448' (Module coreir_reg)
  wire  reg_448__clk;
  wire [15:0] reg_448__in;
  wire [15:0] reg_448__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_448(
    .clk(reg_448__clk),
    .in(reg_448__in),
    .out(reg_448__out)
  );

  //Wire declarations for instance 'reg_449' (Module coreir_reg)
  wire  reg_449__clk;
  wire [15:0] reg_449__in;
  wire [15:0] reg_449__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_449(
    .clk(reg_449__clk),
    .in(reg_449__in),
    .out(reg_449__out)
  );

  //Wire declarations for instance 'reg_45' (Module coreir_reg)
  wire  reg_45__clk;
  wire [15:0] reg_45__in;
  wire [15:0] reg_45__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_45(
    .clk(reg_45__clk),
    .in(reg_45__in),
    .out(reg_45__out)
  );

  //Wire declarations for instance 'reg_450' (Module coreir_reg)
  wire  reg_450__clk;
  wire [15:0] reg_450__in;
  wire [15:0] reg_450__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_450(
    .clk(reg_450__clk),
    .in(reg_450__in),
    .out(reg_450__out)
  );

  //Wire declarations for instance 'reg_451' (Module coreir_reg)
  wire  reg_451__clk;
  wire [15:0] reg_451__in;
  wire [15:0] reg_451__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_451(
    .clk(reg_451__clk),
    .in(reg_451__in),
    .out(reg_451__out)
  );

  //Wire declarations for instance 'reg_452' (Module coreir_reg)
  wire  reg_452__clk;
  wire [15:0] reg_452__in;
  wire [15:0] reg_452__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_452(
    .clk(reg_452__clk),
    .in(reg_452__in),
    .out(reg_452__out)
  );

  //Wire declarations for instance 'reg_453' (Module coreir_reg)
  wire  reg_453__clk;
  wire [15:0] reg_453__in;
  wire [15:0] reg_453__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_453(
    .clk(reg_453__clk),
    .in(reg_453__in),
    .out(reg_453__out)
  );

  //Wire declarations for instance 'reg_454' (Module coreir_reg)
  wire  reg_454__clk;
  wire [15:0] reg_454__in;
  wire [15:0] reg_454__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_454(
    .clk(reg_454__clk),
    .in(reg_454__in),
    .out(reg_454__out)
  );

  //Wire declarations for instance 'reg_455' (Module coreir_reg)
  wire  reg_455__clk;
  wire [15:0] reg_455__in;
  wire [15:0] reg_455__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_455(
    .clk(reg_455__clk),
    .in(reg_455__in),
    .out(reg_455__out)
  );

  //Wire declarations for instance 'reg_456' (Module coreir_reg)
  wire  reg_456__clk;
  wire [15:0] reg_456__in;
  wire [15:0] reg_456__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_456(
    .clk(reg_456__clk),
    .in(reg_456__in),
    .out(reg_456__out)
  );

  //Wire declarations for instance 'reg_457' (Module coreir_reg)
  wire  reg_457__clk;
  wire [15:0] reg_457__in;
  wire [15:0] reg_457__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_457(
    .clk(reg_457__clk),
    .in(reg_457__in),
    .out(reg_457__out)
  );

  //Wire declarations for instance 'reg_458' (Module coreir_reg)
  wire  reg_458__clk;
  wire [15:0] reg_458__in;
  wire [15:0] reg_458__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_458(
    .clk(reg_458__clk),
    .in(reg_458__in),
    .out(reg_458__out)
  );

  //Wire declarations for instance 'reg_459' (Module coreir_reg)
  wire  reg_459__clk;
  wire [15:0] reg_459__in;
  wire [15:0] reg_459__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_459(
    .clk(reg_459__clk),
    .in(reg_459__in),
    .out(reg_459__out)
  );

  //Wire declarations for instance 'reg_46' (Module coreir_reg)
  wire  reg_46__clk;
  wire [15:0] reg_46__in;
  wire [15:0] reg_46__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_46(
    .clk(reg_46__clk),
    .in(reg_46__in),
    .out(reg_46__out)
  );

  //Wire declarations for instance 'reg_460' (Module coreir_reg)
  wire  reg_460__clk;
  wire [15:0] reg_460__in;
  wire [15:0] reg_460__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_460(
    .clk(reg_460__clk),
    .in(reg_460__in),
    .out(reg_460__out)
  );

  //Wire declarations for instance 'reg_461' (Module coreir_reg)
  wire  reg_461__clk;
  wire [15:0] reg_461__in;
  wire [15:0] reg_461__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_461(
    .clk(reg_461__clk),
    .in(reg_461__in),
    .out(reg_461__out)
  );

  //Wire declarations for instance 'reg_462' (Module coreir_reg)
  wire  reg_462__clk;
  wire [15:0] reg_462__in;
  wire [15:0] reg_462__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_462(
    .clk(reg_462__clk),
    .in(reg_462__in),
    .out(reg_462__out)
  );

  //Wire declarations for instance 'reg_463' (Module coreir_reg)
  wire  reg_463__clk;
  wire [15:0] reg_463__in;
  wire [15:0] reg_463__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_463(
    .clk(reg_463__clk),
    .in(reg_463__in),
    .out(reg_463__out)
  );

  //Wire declarations for instance 'reg_464' (Module coreir_reg)
  wire  reg_464__clk;
  wire [15:0] reg_464__in;
  wire [15:0] reg_464__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_464(
    .clk(reg_464__clk),
    .in(reg_464__in),
    .out(reg_464__out)
  );

  //Wire declarations for instance 'reg_465' (Module coreir_reg)
  wire  reg_465__clk;
  wire [15:0] reg_465__in;
  wire [15:0] reg_465__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_465(
    .clk(reg_465__clk),
    .in(reg_465__in),
    .out(reg_465__out)
  );

  //Wire declarations for instance 'reg_466' (Module coreir_reg)
  wire  reg_466__clk;
  wire [15:0] reg_466__in;
  wire [15:0] reg_466__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_466(
    .clk(reg_466__clk),
    .in(reg_466__in),
    .out(reg_466__out)
  );

  //Wire declarations for instance 'reg_467' (Module coreir_reg)
  wire  reg_467__clk;
  wire [15:0] reg_467__in;
  wire [15:0] reg_467__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_467(
    .clk(reg_467__clk),
    .in(reg_467__in),
    .out(reg_467__out)
  );

  //Wire declarations for instance 'reg_468' (Module coreir_reg)
  wire  reg_468__clk;
  wire [15:0] reg_468__in;
  wire [15:0] reg_468__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_468(
    .clk(reg_468__clk),
    .in(reg_468__in),
    .out(reg_468__out)
  );

  //Wire declarations for instance 'reg_469' (Module coreir_reg)
  wire  reg_469__clk;
  wire [15:0] reg_469__in;
  wire [15:0] reg_469__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_469(
    .clk(reg_469__clk),
    .in(reg_469__in),
    .out(reg_469__out)
  );

  //Wire declarations for instance 'reg_47' (Module coreir_reg)
  wire  reg_47__clk;
  wire [15:0] reg_47__in;
  wire [15:0] reg_47__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_47(
    .clk(reg_47__clk),
    .in(reg_47__in),
    .out(reg_47__out)
  );

  //Wire declarations for instance 'reg_470' (Module coreir_reg)
  wire  reg_470__clk;
  wire [15:0] reg_470__in;
  wire [15:0] reg_470__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_470(
    .clk(reg_470__clk),
    .in(reg_470__in),
    .out(reg_470__out)
  );

  //Wire declarations for instance 'reg_471' (Module coreir_reg)
  wire  reg_471__clk;
  wire [15:0] reg_471__in;
  wire [15:0] reg_471__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_471(
    .clk(reg_471__clk),
    .in(reg_471__in),
    .out(reg_471__out)
  );

  //Wire declarations for instance 'reg_472' (Module coreir_reg)
  wire  reg_472__clk;
  wire [15:0] reg_472__in;
  wire [15:0] reg_472__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_472(
    .clk(reg_472__clk),
    .in(reg_472__in),
    .out(reg_472__out)
  );

  //Wire declarations for instance 'reg_473' (Module coreir_reg)
  wire  reg_473__clk;
  wire [15:0] reg_473__in;
  wire [15:0] reg_473__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_473(
    .clk(reg_473__clk),
    .in(reg_473__in),
    .out(reg_473__out)
  );

  //Wire declarations for instance 'reg_474' (Module coreir_reg)
  wire  reg_474__clk;
  wire [15:0] reg_474__in;
  wire [15:0] reg_474__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_474(
    .clk(reg_474__clk),
    .in(reg_474__in),
    .out(reg_474__out)
  );

  //Wire declarations for instance 'reg_475' (Module coreir_reg)
  wire  reg_475__clk;
  wire [15:0] reg_475__in;
  wire [15:0] reg_475__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_475(
    .clk(reg_475__clk),
    .in(reg_475__in),
    .out(reg_475__out)
  );

  //Wire declarations for instance 'reg_476' (Module coreir_reg)
  wire  reg_476__clk;
  wire [15:0] reg_476__in;
  wire [15:0] reg_476__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_476(
    .clk(reg_476__clk),
    .in(reg_476__in),
    .out(reg_476__out)
  );

  //Wire declarations for instance 'reg_477' (Module coreir_reg)
  wire  reg_477__clk;
  wire [15:0] reg_477__in;
  wire [15:0] reg_477__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_477(
    .clk(reg_477__clk),
    .in(reg_477__in),
    .out(reg_477__out)
  );

  //Wire declarations for instance 'reg_478' (Module coreir_reg)
  wire  reg_478__clk;
  wire [15:0] reg_478__in;
  wire [15:0] reg_478__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_478(
    .clk(reg_478__clk),
    .in(reg_478__in),
    .out(reg_478__out)
  );

  //Wire declarations for instance 'reg_479' (Module coreir_reg)
  wire  reg_479__clk;
  wire [15:0] reg_479__in;
  wire [15:0] reg_479__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_479(
    .clk(reg_479__clk),
    .in(reg_479__in),
    .out(reg_479__out)
  );

  //Wire declarations for instance 'reg_48' (Module coreir_reg)
  wire  reg_48__clk;
  wire [15:0] reg_48__in;
  wire [15:0] reg_48__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_48(
    .clk(reg_48__clk),
    .in(reg_48__in),
    .out(reg_48__out)
  );

  //Wire declarations for instance 'reg_480' (Module coreir_reg)
  wire  reg_480__clk;
  wire [15:0] reg_480__in;
  wire [15:0] reg_480__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_480(
    .clk(reg_480__clk),
    .in(reg_480__in),
    .out(reg_480__out)
  );

  //Wire declarations for instance 'reg_481' (Module coreir_reg)
  wire  reg_481__clk;
  wire [15:0] reg_481__in;
  wire [15:0] reg_481__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_481(
    .clk(reg_481__clk),
    .in(reg_481__in),
    .out(reg_481__out)
  );

  //Wire declarations for instance 'reg_482' (Module coreir_reg)
  wire  reg_482__clk;
  wire [15:0] reg_482__in;
  wire [15:0] reg_482__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_482(
    .clk(reg_482__clk),
    .in(reg_482__in),
    .out(reg_482__out)
  );

  //Wire declarations for instance 'reg_483' (Module coreir_reg)
  wire  reg_483__clk;
  wire [15:0] reg_483__in;
  wire [15:0] reg_483__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_483(
    .clk(reg_483__clk),
    .in(reg_483__in),
    .out(reg_483__out)
  );

  //Wire declarations for instance 'reg_484' (Module coreir_reg)
  wire  reg_484__clk;
  wire [15:0] reg_484__in;
  wire [15:0] reg_484__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_484(
    .clk(reg_484__clk),
    .in(reg_484__in),
    .out(reg_484__out)
  );

  //Wire declarations for instance 'reg_485' (Module coreir_reg)
  wire  reg_485__clk;
  wire [15:0] reg_485__in;
  wire [15:0] reg_485__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_485(
    .clk(reg_485__clk),
    .in(reg_485__in),
    .out(reg_485__out)
  );

  //Wire declarations for instance 'reg_486' (Module coreir_reg)
  wire  reg_486__clk;
  wire [15:0] reg_486__in;
  wire [15:0] reg_486__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_486(
    .clk(reg_486__clk),
    .in(reg_486__in),
    .out(reg_486__out)
  );

  //Wire declarations for instance 'reg_487' (Module coreir_reg)
  wire  reg_487__clk;
  wire [15:0] reg_487__in;
  wire [15:0] reg_487__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_487(
    .clk(reg_487__clk),
    .in(reg_487__in),
    .out(reg_487__out)
  );

  //Wire declarations for instance 'reg_488' (Module coreir_reg)
  wire  reg_488__clk;
  wire [15:0] reg_488__in;
  wire [15:0] reg_488__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_488(
    .clk(reg_488__clk),
    .in(reg_488__in),
    .out(reg_488__out)
  );

  //Wire declarations for instance 'reg_489' (Module coreir_reg)
  wire  reg_489__clk;
  wire [15:0] reg_489__in;
  wire [15:0] reg_489__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_489(
    .clk(reg_489__clk),
    .in(reg_489__in),
    .out(reg_489__out)
  );

  //Wire declarations for instance 'reg_49' (Module coreir_reg)
  wire  reg_49__clk;
  wire [15:0] reg_49__in;
  wire [15:0] reg_49__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_49(
    .clk(reg_49__clk),
    .in(reg_49__in),
    .out(reg_49__out)
  );

  //Wire declarations for instance 'reg_490' (Module coreir_reg)
  wire  reg_490__clk;
  wire [15:0] reg_490__in;
  wire [15:0] reg_490__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_490(
    .clk(reg_490__clk),
    .in(reg_490__in),
    .out(reg_490__out)
  );

  //Wire declarations for instance 'reg_491' (Module coreir_reg)
  wire  reg_491__clk;
  wire [15:0] reg_491__in;
  wire [15:0] reg_491__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_491(
    .clk(reg_491__clk),
    .in(reg_491__in),
    .out(reg_491__out)
  );

  //Wire declarations for instance 'reg_492' (Module coreir_reg)
  wire  reg_492__clk;
  wire [15:0] reg_492__in;
  wire [15:0] reg_492__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_492(
    .clk(reg_492__clk),
    .in(reg_492__in),
    .out(reg_492__out)
  );

  //Wire declarations for instance 'reg_493' (Module coreir_reg)
  wire  reg_493__clk;
  wire [15:0] reg_493__in;
  wire [15:0] reg_493__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_493(
    .clk(reg_493__clk),
    .in(reg_493__in),
    .out(reg_493__out)
  );

  //Wire declarations for instance 'reg_494' (Module coreir_reg)
  wire  reg_494__clk;
  wire [15:0] reg_494__in;
  wire [15:0] reg_494__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_494(
    .clk(reg_494__clk),
    .in(reg_494__in),
    .out(reg_494__out)
  );

  //Wire declarations for instance 'reg_495' (Module coreir_reg)
  wire  reg_495__clk;
  wire [15:0] reg_495__in;
  wire [15:0] reg_495__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_495(
    .clk(reg_495__clk),
    .in(reg_495__in),
    .out(reg_495__out)
  );

  //Wire declarations for instance 'reg_496' (Module coreir_reg)
  wire  reg_496__clk;
  wire [15:0] reg_496__in;
  wire [15:0] reg_496__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_496(
    .clk(reg_496__clk),
    .in(reg_496__in),
    .out(reg_496__out)
  );

  //Wire declarations for instance 'reg_497' (Module coreir_reg)
  wire  reg_497__clk;
  wire [15:0] reg_497__in;
  wire [15:0] reg_497__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_497(
    .clk(reg_497__clk),
    .in(reg_497__in),
    .out(reg_497__out)
  );

  //Wire declarations for instance 'reg_498' (Module coreir_reg)
  wire  reg_498__clk;
  wire [15:0] reg_498__in;
  wire [15:0] reg_498__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_498(
    .clk(reg_498__clk),
    .in(reg_498__in),
    .out(reg_498__out)
  );

  //Wire declarations for instance 'reg_499' (Module coreir_reg)
  wire  reg_499__clk;
  wire [15:0] reg_499__in;
  wire [15:0] reg_499__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_499(
    .clk(reg_499__clk),
    .in(reg_499__in),
    .out(reg_499__out)
  );

  //Wire declarations for instance 'reg_5' (Module coreir_reg)
  wire  reg_5__clk;
  wire [15:0] reg_5__in;
  wire [15:0] reg_5__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_5(
    .clk(reg_5__clk),
    .in(reg_5__in),
    .out(reg_5__out)
  );

  //Wire declarations for instance 'reg_50' (Module coreir_reg)
  wire  reg_50__clk;
  wire [15:0] reg_50__in;
  wire [15:0] reg_50__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_50(
    .clk(reg_50__clk),
    .in(reg_50__in),
    .out(reg_50__out)
  );

  //Wire declarations for instance 'reg_500' (Module coreir_reg)
  wire  reg_500__clk;
  wire [15:0] reg_500__in;
  wire [15:0] reg_500__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_500(
    .clk(reg_500__clk),
    .in(reg_500__in),
    .out(reg_500__out)
  );

  //Wire declarations for instance 'reg_501' (Module coreir_reg)
  wire  reg_501__clk;
  wire [15:0] reg_501__in;
  wire [15:0] reg_501__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_501(
    .clk(reg_501__clk),
    .in(reg_501__in),
    .out(reg_501__out)
  );

  //Wire declarations for instance 'reg_502' (Module coreir_reg)
  wire  reg_502__clk;
  wire [15:0] reg_502__in;
  wire [15:0] reg_502__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_502(
    .clk(reg_502__clk),
    .in(reg_502__in),
    .out(reg_502__out)
  );

  //Wire declarations for instance 'reg_503' (Module coreir_reg)
  wire  reg_503__clk;
  wire [15:0] reg_503__in;
  wire [15:0] reg_503__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_503(
    .clk(reg_503__clk),
    .in(reg_503__in),
    .out(reg_503__out)
  );

  //Wire declarations for instance 'reg_504' (Module coreir_reg)
  wire  reg_504__clk;
  wire [15:0] reg_504__in;
  wire [15:0] reg_504__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_504(
    .clk(reg_504__clk),
    .in(reg_504__in),
    .out(reg_504__out)
  );

  //Wire declarations for instance 'reg_505' (Module coreir_reg)
  wire  reg_505__clk;
  wire [15:0] reg_505__in;
  wire [15:0] reg_505__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_505(
    .clk(reg_505__clk),
    .in(reg_505__in),
    .out(reg_505__out)
  );

  //Wire declarations for instance 'reg_506' (Module coreir_reg)
  wire  reg_506__clk;
  wire [15:0] reg_506__in;
  wire [15:0] reg_506__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_506(
    .clk(reg_506__clk),
    .in(reg_506__in),
    .out(reg_506__out)
  );

  //Wire declarations for instance 'reg_507' (Module coreir_reg)
  wire  reg_507__clk;
  wire [15:0] reg_507__in;
  wire [15:0] reg_507__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_507(
    .clk(reg_507__clk),
    .in(reg_507__in),
    .out(reg_507__out)
  );

  //Wire declarations for instance 'reg_508' (Module coreir_reg)
  wire  reg_508__clk;
  wire [15:0] reg_508__in;
  wire [15:0] reg_508__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_508(
    .clk(reg_508__clk),
    .in(reg_508__in),
    .out(reg_508__out)
  );

  //Wire declarations for instance 'reg_509' (Module coreir_reg)
  wire  reg_509__clk;
  wire [15:0] reg_509__in;
  wire [15:0] reg_509__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_509(
    .clk(reg_509__clk),
    .in(reg_509__in),
    .out(reg_509__out)
  );

  //Wire declarations for instance 'reg_51' (Module coreir_reg)
  wire  reg_51__clk;
  wire [15:0] reg_51__in;
  wire [15:0] reg_51__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_51(
    .clk(reg_51__clk),
    .in(reg_51__in),
    .out(reg_51__out)
  );

  //Wire declarations for instance 'reg_510' (Module coreir_reg)
  wire  reg_510__clk;
  wire [15:0] reg_510__in;
  wire [15:0] reg_510__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_510(
    .clk(reg_510__clk),
    .in(reg_510__in),
    .out(reg_510__out)
  );

  //Wire declarations for instance 'reg_511' (Module coreir_reg)
  wire  reg_511__clk;
  wire [15:0] reg_511__in;
  wire [15:0] reg_511__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_511(
    .clk(reg_511__clk),
    .in(reg_511__in),
    .out(reg_511__out)
  );

  //Wire declarations for instance 'reg_512' (Module coreir_reg)
  wire  reg_512__clk;
  wire [15:0] reg_512__in;
  wire [15:0] reg_512__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_512(
    .clk(reg_512__clk),
    .in(reg_512__in),
    .out(reg_512__out)
  );

  //Wire declarations for instance 'reg_513' (Module coreir_reg)
  wire  reg_513__clk;
  wire [15:0] reg_513__in;
  wire [15:0] reg_513__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_513(
    .clk(reg_513__clk),
    .in(reg_513__in),
    .out(reg_513__out)
  );

  //Wire declarations for instance 'reg_514' (Module coreir_reg)
  wire  reg_514__clk;
  wire [15:0] reg_514__in;
  wire [15:0] reg_514__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_514(
    .clk(reg_514__clk),
    .in(reg_514__in),
    .out(reg_514__out)
  );

  //Wire declarations for instance 'reg_515' (Module coreir_reg)
  wire  reg_515__clk;
  wire [15:0] reg_515__in;
  wire [15:0] reg_515__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_515(
    .clk(reg_515__clk),
    .in(reg_515__in),
    .out(reg_515__out)
  );

  //Wire declarations for instance 'reg_516' (Module coreir_reg)
  wire  reg_516__clk;
  wire [15:0] reg_516__in;
  wire [15:0] reg_516__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_516(
    .clk(reg_516__clk),
    .in(reg_516__in),
    .out(reg_516__out)
  );

  //Wire declarations for instance 'reg_517' (Module coreir_reg)
  wire  reg_517__clk;
  wire [15:0] reg_517__in;
  wire [15:0] reg_517__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_517(
    .clk(reg_517__clk),
    .in(reg_517__in),
    .out(reg_517__out)
  );

  //Wire declarations for instance 'reg_518' (Module coreir_reg)
  wire  reg_518__clk;
  wire [15:0] reg_518__in;
  wire [15:0] reg_518__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_518(
    .clk(reg_518__clk),
    .in(reg_518__in),
    .out(reg_518__out)
  );

  //Wire declarations for instance 'reg_519' (Module coreir_reg)
  wire  reg_519__clk;
  wire [15:0] reg_519__in;
  wire [15:0] reg_519__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_519(
    .clk(reg_519__clk),
    .in(reg_519__in),
    .out(reg_519__out)
  );

  //Wire declarations for instance 'reg_52' (Module coreir_reg)
  wire  reg_52__clk;
  wire [15:0] reg_52__in;
  wire [15:0] reg_52__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_52(
    .clk(reg_52__clk),
    .in(reg_52__in),
    .out(reg_52__out)
  );

  //Wire declarations for instance 'reg_520' (Module coreir_reg)
  wire  reg_520__clk;
  wire [15:0] reg_520__in;
  wire [15:0] reg_520__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_520(
    .clk(reg_520__clk),
    .in(reg_520__in),
    .out(reg_520__out)
  );

  //Wire declarations for instance 'reg_521' (Module coreir_reg)
  wire  reg_521__clk;
  wire [15:0] reg_521__in;
  wire [15:0] reg_521__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_521(
    .clk(reg_521__clk),
    .in(reg_521__in),
    .out(reg_521__out)
  );

  //Wire declarations for instance 'reg_522' (Module coreir_reg)
  wire  reg_522__clk;
  wire [15:0] reg_522__in;
  wire [15:0] reg_522__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_522(
    .clk(reg_522__clk),
    .in(reg_522__in),
    .out(reg_522__out)
  );

  //Wire declarations for instance 'reg_523' (Module coreir_reg)
  wire  reg_523__clk;
  wire [15:0] reg_523__in;
  wire [15:0] reg_523__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_523(
    .clk(reg_523__clk),
    .in(reg_523__in),
    .out(reg_523__out)
  );

  //Wire declarations for instance 'reg_524' (Module coreir_reg)
  wire  reg_524__clk;
  wire [15:0] reg_524__in;
  wire [15:0] reg_524__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_524(
    .clk(reg_524__clk),
    .in(reg_524__in),
    .out(reg_524__out)
  );

  //Wire declarations for instance 'reg_525' (Module coreir_reg)
  wire  reg_525__clk;
  wire [15:0] reg_525__in;
  wire [15:0] reg_525__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_525(
    .clk(reg_525__clk),
    .in(reg_525__in),
    .out(reg_525__out)
  );

  //Wire declarations for instance 'reg_526' (Module coreir_reg)
  wire  reg_526__clk;
  wire [15:0] reg_526__in;
  wire [15:0] reg_526__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_526(
    .clk(reg_526__clk),
    .in(reg_526__in),
    .out(reg_526__out)
  );

  //Wire declarations for instance 'reg_527' (Module coreir_reg)
  wire  reg_527__clk;
  wire [15:0] reg_527__in;
  wire [15:0] reg_527__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_527(
    .clk(reg_527__clk),
    .in(reg_527__in),
    .out(reg_527__out)
  );

  //Wire declarations for instance 'reg_528' (Module coreir_reg)
  wire  reg_528__clk;
  wire [15:0] reg_528__in;
  wire [15:0] reg_528__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_528(
    .clk(reg_528__clk),
    .in(reg_528__in),
    .out(reg_528__out)
  );

  //Wire declarations for instance 'reg_529' (Module coreir_reg)
  wire  reg_529__clk;
  wire [15:0] reg_529__in;
  wire [15:0] reg_529__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_529(
    .clk(reg_529__clk),
    .in(reg_529__in),
    .out(reg_529__out)
  );

  //Wire declarations for instance 'reg_53' (Module coreir_reg)
  wire  reg_53__clk;
  wire [15:0] reg_53__in;
  wire [15:0] reg_53__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_53(
    .clk(reg_53__clk),
    .in(reg_53__in),
    .out(reg_53__out)
  );

  //Wire declarations for instance 'reg_530' (Module coreir_reg)
  wire  reg_530__clk;
  wire [15:0] reg_530__in;
  wire [15:0] reg_530__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_530(
    .clk(reg_530__clk),
    .in(reg_530__in),
    .out(reg_530__out)
  );

  //Wire declarations for instance 'reg_531' (Module coreir_reg)
  wire  reg_531__clk;
  wire [15:0] reg_531__in;
  wire [15:0] reg_531__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_531(
    .clk(reg_531__clk),
    .in(reg_531__in),
    .out(reg_531__out)
  );

  //Wire declarations for instance 'reg_532' (Module coreir_reg)
  wire  reg_532__clk;
  wire [15:0] reg_532__in;
  wire [15:0] reg_532__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_532(
    .clk(reg_532__clk),
    .in(reg_532__in),
    .out(reg_532__out)
  );

  //Wire declarations for instance 'reg_533' (Module coreir_reg)
  wire  reg_533__clk;
  wire [15:0] reg_533__in;
  wire [15:0] reg_533__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_533(
    .clk(reg_533__clk),
    .in(reg_533__in),
    .out(reg_533__out)
  );

  //Wire declarations for instance 'reg_534' (Module coreir_reg)
  wire  reg_534__clk;
  wire [15:0] reg_534__in;
  wire [15:0] reg_534__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_534(
    .clk(reg_534__clk),
    .in(reg_534__in),
    .out(reg_534__out)
  );

  //Wire declarations for instance 'reg_535' (Module coreir_reg)
  wire  reg_535__clk;
  wire [15:0] reg_535__in;
  wire [15:0] reg_535__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_535(
    .clk(reg_535__clk),
    .in(reg_535__in),
    .out(reg_535__out)
  );

  //Wire declarations for instance 'reg_536' (Module coreir_reg)
  wire  reg_536__clk;
  wire [15:0] reg_536__in;
  wire [15:0] reg_536__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_536(
    .clk(reg_536__clk),
    .in(reg_536__in),
    .out(reg_536__out)
  );

  //Wire declarations for instance 'reg_537' (Module coreir_reg)
  wire  reg_537__clk;
  wire [15:0] reg_537__in;
  wire [15:0] reg_537__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_537(
    .clk(reg_537__clk),
    .in(reg_537__in),
    .out(reg_537__out)
  );

  //Wire declarations for instance 'reg_538' (Module coreir_reg)
  wire  reg_538__clk;
  wire [15:0] reg_538__in;
  wire [15:0] reg_538__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_538(
    .clk(reg_538__clk),
    .in(reg_538__in),
    .out(reg_538__out)
  );

  //Wire declarations for instance 'reg_539' (Module coreir_reg)
  wire  reg_539__clk;
  wire [15:0] reg_539__in;
  wire [15:0] reg_539__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_539(
    .clk(reg_539__clk),
    .in(reg_539__in),
    .out(reg_539__out)
  );

  //Wire declarations for instance 'reg_54' (Module coreir_reg)
  wire  reg_54__clk;
  wire [15:0] reg_54__in;
  wire [15:0] reg_54__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_54(
    .clk(reg_54__clk),
    .in(reg_54__in),
    .out(reg_54__out)
  );

  //Wire declarations for instance 'reg_540' (Module coreir_reg)
  wire  reg_540__clk;
  wire [15:0] reg_540__in;
  wire [15:0] reg_540__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_540(
    .clk(reg_540__clk),
    .in(reg_540__in),
    .out(reg_540__out)
  );

  //Wire declarations for instance 'reg_541' (Module coreir_reg)
  wire  reg_541__clk;
  wire [15:0] reg_541__in;
  wire [15:0] reg_541__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_541(
    .clk(reg_541__clk),
    .in(reg_541__in),
    .out(reg_541__out)
  );

  //Wire declarations for instance 'reg_542' (Module coreir_reg)
  wire  reg_542__clk;
  wire [15:0] reg_542__in;
  wire [15:0] reg_542__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_542(
    .clk(reg_542__clk),
    .in(reg_542__in),
    .out(reg_542__out)
  );

  //Wire declarations for instance 'reg_543' (Module coreir_reg)
  wire  reg_543__clk;
  wire [15:0] reg_543__in;
  wire [15:0] reg_543__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_543(
    .clk(reg_543__clk),
    .in(reg_543__in),
    .out(reg_543__out)
  );

  //Wire declarations for instance 'reg_544' (Module coreir_reg)
  wire  reg_544__clk;
  wire [15:0] reg_544__in;
  wire [15:0] reg_544__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_544(
    .clk(reg_544__clk),
    .in(reg_544__in),
    .out(reg_544__out)
  );

  //Wire declarations for instance 'reg_545' (Module coreir_reg)
  wire  reg_545__clk;
  wire [15:0] reg_545__in;
  wire [15:0] reg_545__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_545(
    .clk(reg_545__clk),
    .in(reg_545__in),
    .out(reg_545__out)
  );

  //Wire declarations for instance 'reg_546' (Module coreir_reg)
  wire  reg_546__clk;
  wire [15:0] reg_546__in;
  wire [15:0] reg_546__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_546(
    .clk(reg_546__clk),
    .in(reg_546__in),
    .out(reg_546__out)
  );

  //Wire declarations for instance 'reg_547' (Module coreir_reg)
  wire  reg_547__clk;
  wire [15:0] reg_547__in;
  wire [15:0] reg_547__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_547(
    .clk(reg_547__clk),
    .in(reg_547__in),
    .out(reg_547__out)
  );

  //Wire declarations for instance 'reg_548' (Module coreir_reg)
  wire  reg_548__clk;
  wire [15:0] reg_548__in;
  wire [15:0] reg_548__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_548(
    .clk(reg_548__clk),
    .in(reg_548__in),
    .out(reg_548__out)
  );

  //Wire declarations for instance 'reg_549' (Module coreir_reg)
  wire  reg_549__clk;
  wire [15:0] reg_549__in;
  wire [15:0] reg_549__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_549(
    .clk(reg_549__clk),
    .in(reg_549__in),
    .out(reg_549__out)
  );

  //Wire declarations for instance 'reg_55' (Module coreir_reg)
  wire  reg_55__clk;
  wire [15:0] reg_55__in;
  wire [15:0] reg_55__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_55(
    .clk(reg_55__clk),
    .in(reg_55__in),
    .out(reg_55__out)
  );

  //Wire declarations for instance 'reg_550' (Module coreir_reg)
  wire  reg_550__clk;
  wire [15:0] reg_550__in;
  wire [15:0] reg_550__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_550(
    .clk(reg_550__clk),
    .in(reg_550__in),
    .out(reg_550__out)
  );

  //Wire declarations for instance 'reg_551' (Module coreir_reg)
  wire  reg_551__clk;
  wire [15:0] reg_551__in;
  wire [15:0] reg_551__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_551(
    .clk(reg_551__clk),
    .in(reg_551__in),
    .out(reg_551__out)
  );

  //Wire declarations for instance 'reg_552' (Module coreir_reg)
  wire  reg_552__clk;
  wire [15:0] reg_552__in;
  wire [15:0] reg_552__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_552(
    .clk(reg_552__clk),
    .in(reg_552__in),
    .out(reg_552__out)
  );

  //Wire declarations for instance 'reg_553' (Module coreir_reg)
  wire  reg_553__clk;
  wire [15:0] reg_553__in;
  wire [15:0] reg_553__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_553(
    .clk(reg_553__clk),
    .in(reg_553__in),
    .out(reg_553__out)
  );

  //Wire declarations for instance 'reg_554' (Module coreir_reg)
  wire  reg_554__clk;
  wire [15:0] reg_554__in;
  wire [15:0] reg_554__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_554(
    .clk(reg_554__clk),
    .in(reg_554__in),
    .out(reg_554__out)
  );

  //Wire declarations for instance 'reg_555' (Module coreir_reg)
  wire  reg_555__clk;
  wire [15:0] reg_555__in;
  wire [15:0] reg_555__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_555(
    .clk(reg_555__clk),
    .in(reg_555__in),
    .out(reg_555__out)
  );

  //Wire declarations for instance 'reg_556' (Module coreir_reg)
  wire  reg_556__clk;
  wire [15:0] reg_556__in;
  wire [15:0] reg_556__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_556(
    .clk(reg_556__clk),
    .in(reg_556__in),
    .out(reg_556__out)
  );

  //Wire declarations for instance 'reg_557' (Module coreir_reg)
  wire  reg_557__clk;
  wire [15:0] reg_557__in;
  wire [15:0] reg_557__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_557(
    .clk(reg_557__clk),
    .in(reg_557__in),
    .out(reg_557__out)
  );

  //Wire declarations for instance 'reg_558' (Module coreir_reg)
  wire  reg_558__clk;
  wire [15:0] reg_558__in;
  wire [15:0] reg_558__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_558(
    .clk(reg_558__clk),
    .in(reg_558__in),
    .out(reg_558__out)
  );

  //Wire declarations for instance 'reg_559' (Module coreir_reg)
  wire  reg_559__clk;
  wire [15:0] reg_559__in;
  wire [15:0] reg_559__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_559(
    .clk(reg_559__clk),
    .in(reg_559__in),
    .out(reg_559__out)
  );

  //Wire declarations for instance 'reg_56' (Module coreir_reg)
  wire  reg_56__clk;
  wire [15:0] reg_56__in;
  wire [15:0] reg_56__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_56(
    .clk(reg_56__clk),
    .in(reg_56__in),
    .out(reg_56__out)
  );

  //Wire declarations for instance 'reg_560' (Module coreir_reg)
  wire  reg_560__clk;
  wire [15:0] reg_560__in;
  wire [15:0] reg_560__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_560(
    .clk(reg_560__clk),
    .in(reg_560__in),
    .out(reg_560__out)
  );

  //Wire declarations for instance 'reg_561' (Module coreir_reg)
  wire  reg_561__clk;
  wire [15:0] reg_561__in;
  wire [15:0] reg_561__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_561(
    .clk(reg_561__clk),
    .in(reg_561__in),
    .out(reg_561__out)
  );

  //Wire declarations for instance 'reg_562' (Module coreir_reg)
  wire  reg_562__clk;
  wire [15:0] reg_562__in;
  wire [15:0] reg_562__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_562(
    .clk(reg_562__clk),
    .in(reg_562__in),
    .out(reg_562__out)
  );

  //Wire declarations for instance 'reg_563' (Module coreir_reg)
  wire  reg_563__clk;
  wire [15:0] reg_563__in;
  wire [15:0] reg_563__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_563(
    .clk(reg_563__clk),
    .in(reg_563__in),
    .out(reg_563__out)
  );

  //Wire declarations for instance 'reg_564' (Module coreir_reg)
  wire  reg_564__clk;
  wire [15:0] reg_564__in;
  wire [15:0] reg_564__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_564(
    .clk(reg_564__clk),
    .in(reg_564__in),
    .out(reg_564__out)
  );

  //Wire declarations for instance 'reg_565' (Module coreir_reg)
  wire  reg_565__clk;
  wire [15:0] reg_565__in;
  wire [15:0] reg_565__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_565(
    .clk(reg_565__clk),
    .in(reg_565__in),
    .out(reg_565__out)
  );

  //Wire declarations for instance 'reg_566' (Module coreir_reg)
  wire  reg_566__clk;
  wire [15:0] reg_566__in;
  wire [15:0] reg_566__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_566(
    .clk(reg_566__clk),
    .in(reg_566__in),
    .out(reg_566__out)
  );

  //Wire declarations for instance 'reg_567' (Module coreir_reg)
  wire  reg_567__clk;
  wire [15:0] reg_567__in;
  wire [15:0] reg_567__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_567(
    .clk(reg_567__clk),
    .in(reg_567__in),
    .out(reg_567__out)
  );

  //Wire declarations for instance 'reg_568' (Module coreir_reg)
  wire  reg_568__clk;
  wire [15:0] reg_568__in;
  wire [15:0] reg_568__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_568(
    .clk(reg_568__clk),
    .in(reg_568__in),
    .out(reg_568__out)
  );

  //Wire declarations for instance 'reg_569' (Module coreir_reg)
  wire  reg_569__clk;
  wire [15:0] reg_569__in;
  wire [15:0] reg_569__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_569(
    .clk(reg_569__clk),
    .in(reg_569__in),
    .out(reg_569__out)
  );

  //Wire declarations for instance 'reg_57' (Module coreir_reg)
  wire  reg_57__clk;
  wire [15:0] reg_57__in;
  wire [15:0] reg_57__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_57(
    .clk(reg_57__clk),
    .in(reg_57__in),
    .out(reg_57__out)
  );

  //Wire declarations for instance 'reg_570' (Module coreir_reg)
  wire  reg_570__clk;
  wire [15:0] reg_570__in;
  wire [15:0] reg_570__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_570(
    .clk(reg_570__clk),
    .in(reg_570__in),
    .out(reg_570__out)
  );

  //Wire declarations for instance 'reg_571' (Module coreir_reg)
  wire  reg_571__clk;
  wire [15:0] reg_571__in;
  wire [15:0] reg_571__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_571(
    .clk(reg_571__clk),
    .in(reg_571__in),
    .out(reg_571__out)
  );

  //Wire declarations for instance 'reg_572' (Module coreir_reg)
  wire  reg_572__clk;
  wire [15:0] reg_572__in;
  wire [15:0] reg_572__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_572(
    .clk(reg_572__clk),
    .in(reg_572__in),
    .out(reg_572__out)
  );

  //Wire declarations for instance 'reg_573' (Module coreir_reg)
  wire  reg_573__clk;
  wire [15:0] reg_573__in;
  wire [15:0] reg_573__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_573(
    .clk(reg_573__clk),
    .in(reg_573__in),
    .out(reg_573__out)
  );

  //Wire declarations for instance 'reg_574' (Module coreir_reg)
  wire  reg_574__clk;
  wire [15:0] reg_574__in;
  wire [15:0] reg_574__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_574(
    .clk(reg_574__clk),
    .in(reg_574__in),
    .out(reg_574__out)
  );

  //Wire declarations for instance 'reg_575' (Module coreir_reg)
  wire  reg_575__clk;
  wire [15:0] reg_575__in;
  wire [15:0] reg_575__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_575(
    .clk(reg_575__clk),
    .in(reg_575__in),
    .out(reg_575__out)
  );

  //Wire declarations for instance 'reg_576' (Module coreir_reg)
  wire  reg_576__clk;
  wire [15:0] reg_576__in;
  wire [15:0] reg_576__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_576(
    .clk(reg_576__clk),
    .in(reg_576__in),
    .out(reg_576__out)
  );

  //Wire declarations for instance 'reg_577' (Module coreir_reg)
  wire  reg_577__clk;
  wire [15:0] reg_577__in;
  wire [15:0] reg_577__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_577(
    .clk(reg_577__clk),
    .in(reg_577__in),
    .out(reg_577__out)
  );

  //Wire declarations for instance 'reg_578' (Module coreir_reg)
  wire  reg_578__clk;
  wire [15:0] reg_578__in;
  wire [15:0] reg_578__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_578(
    .clk(reg_578__clk),
    .in(reg_578__in),
    .out(reg_578__out)
  );

  //Wire declarations for instance 'reg_579' (Module coreir_reg)
  wire  reg_579__clk;
  wire [15:0] reg_579__in;
  wire [15:0] reg_579__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_579(
    .clk(reg_579__clk),
    .in(reg_579__in),
    .out(reg_579__out)
  );

  //Wire declarations for instance 'reg_58' (Module coreir_reg)
  wire  reg_58__clk;
  wire [15:0] reg_58__in;
  wire [15:0] reg_58__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_58(
    .clk(reg_58__clk),
    .in(reg_58__in),
    .out(reg_58__out)
  );

  //Wire declarations for instance 'reg_580' (Module coreir_reg)
  wire  reg_580__clk;
  wire [15:0] reg_580__in;
  wire [15:0] reg_580__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_580(
    .clk(reg_580__clk),
    .in(reg_580__in),
    .out(reg_580__out)
  );

  //Wire declarations for instance 'reg_581' (Module coreir_reg)
  wire  reg_581__clk;
  wire [15:0] reg_581__in;
  wire [15:0] reg_581__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_581(
    .clk(reg_581__clk),
    .in(reg_581__in),
    .out(reg_581__out)
  );

  //Wire declarations for instance 'reg_582' (Module coreir_reg)
  wire  reg_582__clk;
  wire [15:0] reg_582__in;
  wire [15:0] reg_582__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_582(
    .clk(reg_582__clk),
    .in(reg_582__in),
    .out(reg_582__out)
  );

  //Wire declarations for instance 'reg_583' (Module coreir_reg)
  wire  reg_583__clk;
  wire [15:0] reg_583__in;
  wire [15:0] reg_583__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_583(
    .clk(reg_583__clk),
    .in(reg_583__in),
    .out(reg_583__out)
  );

  //Wire declarations for instance 'reg_584' (Module coreir_reg)
  wire  reg_584__clk;
  wire [15:0] reg_584__in;
  wire [15:0] reg_584__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_584(
    .clk(reg_584__clk),
    .in(reg_584__in),
    .out(reg_584__out)
  );

  //Wire declarations for instance 'reg_585' (Module coreir_reg)
  wire  reg_585__clk;
  wire [15:0] reg_585__in;
  wire [15:0] reg_585__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_585(
    .clk(reg_585__clk),
    .in(reg_585__in),
    .out(reg_585__out)
  );

  //Wire declarations for instance 'reg_586' (Module coreir_reg)
  wire  reg_586__clk;
  wire [15:0] reg_586__in;
  wire [15:0] reg_586__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_586(
    .clk(reg_586__clk),
    .in(reg_586__in),
    .out(reg_586__out)
  );

  //Wire declarations for instance 'reg_587' (Module coreir_reg)
  wire  reg_587__clk;
  wire [15:0] reg_587__in;
  wire [15:0] reg_587__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_587(
    .clk(reg_587__clk),
    .in(reg_587__in),
    .out(reg_587__out)
  );

  //Wire declarations for instance 'reg_588' (Module coreir_reg)
  wire  reg_588__clk;
  wire [15:0] reg_588__in;
  wire [15:0] reg_588__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_588(
    .clk(reg_588__clk),
    .in(reg_588__in),
    .out(reg_588__out)
  );

  //Wire declarations for instance 'reg_589' (Module coreir_reg)
  wire  reg_589__clk;
  wire [15:0] reg_589__in;
  wire [15:0] reg_589__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_589(
    .clk(reg_589__clk),
    .in(reg_589__in),
    .out(reg_589__out)
  );

  //Wire declarations for instance 'reg_59' (Module coreir_reg)
  wire  reg_59__clk;
  wire [15:0] reg_59__in;
  wire [15:0] reg_59__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_59(
    .clk(reg_59__clk),
    .in(reg_59__in),
    .out(reg_59__out)
  );

  //Wire declarations for instance 'reg_590' (Module coreir_reg)
  wire  reg_590__clk;
  wire [15:0] reg_590__in;
  wire [15:0] reg_590__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_590(
    .clk(reg_590__clk),
    .in(reg_590__in),
    .out(reg_590__out)
  );

  //Wire declarations for instance 'reg_591' (Module coreir_reg)
  wire  reg_591__clk;
  wire [15:0] reg_591__in;
  wire [15:0] reg_591__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_591(
    .clk(reg_591__clk),
    .in(reg_591__in),
    .out(reg_591__out)
  );

  //Wire declarations for instance 'reg_592' (Module coreir_reg)
  wire  reg_592__clk;
  wire [15:0] reg_592__in;
  wire [15:0] reg_592__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_592(
    .clk(reg_592__clk),
    .in(reg_592__in),
    .out(reg_592__out)
  );

  //Wire declarations for instance 'reg_593' (Module coreir_reg)
  wire  reg_593__clk;
  wire [15:0] reg_593__in;
  wire [15:0] reg_593__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_593(
    .clk(reg_593__clk),
    .in(reg_593__in),
    .out(reg_593__out)
  );

  //Wire declarations for instance 'reg_594' (Module coreir_reg)
  wire  reg_594__clk;
  wire [15:0] reg_594__in;
  wire [15:0] reg_594__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_594(
    .clk(reg_594__clk),
    .in(reg_594__in),
    .out(reg_594__out)
  );

  //Wire declarations for instance 'reg_595' (Module coreir_reg)
  wire  reg_595__clk;
  wire [15:0] reg_595__in;
  wire [15:0] reg_595__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_595(
    .clk(reg_595__clk),
    .in(reg_595__in),
    .out(reg_595__out)
  );

  //Wire declarations for instance 'reg_596' (Module coreir_reg)
  wire  reg_596__clk;
  wire [15:0] reg_596__in;
  wire [15:0] reg_596__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_596(
    .clk(reg_596__clk),
    .in(reg_596__in),
    .out(reg_596__out)
  );

  //Wire declarations for instance 'reg_597' (Module coreir_reg)
  wire  reg_597__clk;
  wire [15:0] reg_597__in;
  wire [15:0] reg_597__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_597(
    .clk(reg_597__clk),
    .in(reg_597__in),
    .out(reg_597__out)
  );

  //Wire declarations for instance 'reg_598' (Module coreir_reg)
  wire  reg_598__clk;
  wire [15:0] reg_598__in;
  wire [15:0] reg_598__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_598(
    .clk(reg_598__clk),
    .in(reg_598__in),
    .out(reg_598__out)
  );

  //Wire declarations for instance 'reg_599' (Module coreir_reg)
  wire  reg_599__clk;
  wire [15:0] reg_599__in;
  wire [15:0] reg_599__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_599(
    .clk(reg_599__clk),
    .in(reg_599__in),
    .out(reg_599__out)
  );

  //Wire declarations for instance 'reg_6' (Module coreir_reg)
  wire  reg_6__clk;
  wire [15:0] reg_6__in;
  wire [15:0] reg_6__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_6(
    .clk(reg_6__clk),
    .in(reg_6__in),
    .out(reg_6__out)
  );

  //Wire declarations for instance 'reg_60' (Module coreir_reg)
  wire  reg_60__clk;
  wire [15:0] reg_60__in;
  wire [15:0] reg_60__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_60(
    .clk(reg_60__clk),
    .in(reg_60__in),
    .out(reg_60__out)
  );

  //Wire declarations for instance 'reg_600' (Module coreir_reg)
  wire  reg_600__clk;
  wire [15:0] reg_600__in;
  wire [15:0] reg_600__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_600(
    .clk(reg_600__clk),
    .in(reg_600__in),
    .out(reg_600__out)
  );

  //Wire declarations for instance 'reg_601' (Module coreir_reg)
  wire  reg_601__clk;
  wire [15:0] reg_601__in;
  wire [15:0] reg_601__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_601(
    .clk(reg_601__clk),
    .in(reg_601__in),
    .out(reg_601__out)
  );

  //Wire declarations for instance 'reg_602' (Module coreir_reg)
  wire  reg_602__clk;
  wire [15:0] reg_602__in;
  wire [15:0] reg_602__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_602(
    .clk(reg_602__clk),
    .in(reg_602__in),
    .out(reg_602__out)
  );

  //Wire declarations for instance 'reg_603' (Module coreir_reg)
  wire  reg_603__clk;
  wire [15:0] reg_603__in;
  wire [15:0] reg_603__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_603(
    .clk(reg_603__clk),
    .in(reg_603__in),
    .out(reg_603__out)
  );

  //Wire declarations for instance 'reg_604' (Module coreir_reg)
  wire  reg_604__clk;
  wire [15:0] reg_604__in;
  wire [15:0] reg_604__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_604(
    .clk(reg_604__clk),
    .in(reg_604__in),
    .out(reg_604__out)
  );

  //Wire declarations for instance 'reg_605' (Module coreir_reg)
  wire  reg_605__clk;
  wire [15:0] reg_605__in;
  wire [15:0] reg_605__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_605(
    .clk(reg_605__clk),
    .in(reg_605__in),
    .out(reg_605__out)
  );

  //Wire declarations for instance 'reg_606' (Module coreir_reg)
  wire  reg_606__clk;
  wire [15:0] reg_606__in;
  wire [15:0] reg_606__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_606(
    .clk(reg_606__clk),
    .in(reg_606__in),
    .out(reg_606__out)
  );

  //Wire declarations for instance 'reg_607' (Module coreir_reg)
  wire  reg_607__clk;
  wire [15:0] reg_607__in;
  wire [15:0] reg_607__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_607(
    .clk(reg_607__clk),
    .in(reg_607__in),
    .out(reg_607__out)
  );

  //Wire declarations for instance 'reg_608' (Module coreir_reg)
  wire  reg_608__clk;
  wire [15:0] reg_608__in;
  wire [15:0] reg_608__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_608(
    .clk(reg_608__clk),
    .in(reg_608__in),
    .out(reg_608__out)
  );

  //Wire declarations for instance 'reg_609' (Module coreir_reg)
  wire  reg_609__clk;
  wire [15:0] reg_609__in;
  wire [15:0] reg_609__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_609(
    .clk(reg_609__clk),
    .in(reg_609__in),
    .out(reg_609__out)
  );

  //Wire declarations for instance 'reg_61' (Module coreir_reg)
  wire  reg_61__clk;
  wire [15:0] reg_61__in;
  wire [15:0] reg_61__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_61(
    .clk(reg_61__clk),
    .in(reg_61__in),
    .out(reg_61__out)
  );

  //Wire declarations for instance 'reg_610' (Module coreir_reg)
  wire  reg_610__clk;
  wire [15:0] reg_610__in;
  wire [15:0] reg_610__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_610(
    .clk(reg_610__clk),
    .in(reg_610__in),
    .out(reg_610__out)
  );

  //Wire declarations for instance 'reg_611' (Module coreir_reg)
  wire  reg_611__clk;
  wire [15:0] reg_611__in;
  wire [15:0] reg_611__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_611(
    .clk(reg_611__clk),
    .in(reg_611__in),
    .out(reg_611__out)
  );

  //Wire declarations for instance 'reg_612' (Module coreir_reg)
  wire  reg_612__clk;
  wire [15:0] reg_612__in;
  wire [15:0] reg_612__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_612(
    .clk(reg_612__clk),
    .in(reg_612__in),
    .out(reg_612__out)
  );

  //Wire declarations for instance 'reg_613' (Module coreir_reg)
  wire  reg_613__clk;
  wire [15:0] reg_613__in;
  wire [15:0] reg_613__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_613(
    .clk(reg_613__clk),
    .in(reg_613__in),
    .out(reg_613__out)
  );

  //Wire declarations for instance 'reg_614' (Module coreir_reg)
  wire  reg_614__clk;
  wire [15:0] reg_614__in;
  wire [15:0] reg_614__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_614(
    .clk(reg_614__clk),
    .in(reg_614__in),
    .out(reg_614__out)
  );

  //Wire declarations for instance 'reg_615' (Module coreir_reg)
  wire  reg_615__clk;
  wire [15:0] reg_615__in;
  wire [15:0] reg_615__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_615(
    .clk(reg_615__clk),
    .in(reg_615__in),
    .out(reg_615__out)
  );

  //Wire declarations for instance 'reg_616' (Module coreir_reg)
  wire  reg_616__clk;
  wire [15:0] reg_616__in;
  wire [15:0] reg_616__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_616(
    .clk(reg_616__clk),
    .in(reg_616__in),
    .out(reg_616__out)
  );

  //Wire declarations for instance 'reg_617' (Module coreir_reg)
  wire  reg_617__clk;
  wire [15:0] reg_617__in;
  wire [15:0] reg_617__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_617(
    .clk(reg_617__clk),
    .in(reg_617__in),
    .out(reg_617__out)
  );

  //Wire declarations for instance 'reg_618' (Module coreir_reg)
  wire  reg_618__clk;
  wire [15:0] reg_618__in;
  wire [15:0] reg_618__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_618(
    .clk(reg_618__clk),
    .in(reg_618__in),
    .out(reg_618__out)
  );

  //Wire declarations for instance 'reg_619' (Module coreir_reg)
  wire  reg_619__clk;
  wire [15:0] reg_619__in;
  wire [15:0] reg_619__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_619(
    .clk(reg_619__clk),
    .in(reg_619__in),
    .out(reg_619__out)
  );

  //Wire declarations for instance 'reg_62' (Module coreir_reg)
  wire  reg_62__clk;
  wire [15:0] reg_62__in;
  wire [15:0] reg_62__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_62(
    .clk(reg_62__clk),
    .in(reg_62__in),
    .out(reg_62__out)
  );

  //Wire declarations for instance 'reg_620' (Module coreir_reg)
  wire  reg_620__clk;
  wire [15:0] reg_620__in;
  wire [15:0] reg_620__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_620(
    .clk(reg_620__clk),
    .in(reg_620__in),
    .out(reg_620__out)
  );

  //Wire declarations for instance 'reg_621' (Module coreir_reg)
  wire  reg_621__clk;
  wire [15:0] reg_621__in;
  wire [15:0] reg_621__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_621(
    .clk(reg_621__clk),
    .in(reg_621__in),
    .out(reg_621__out)
  );

  //Wire declarations for instance 'reg_622' (Module coreir_reg)
  wire  reg_622__clk;
  wire [15:0] reg_622__in;
  wire [15:0] reg_622__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_622(
    .clk(reg_622__clk),
    .in(reg_622__in),
    .out(reg_622__out)
  );

  //Wire declarations for instance 'reg_623' (Module coreir_reg)
  wire  reg_623__clk;
  wire [15:0] reg_623__in;
  wire [15:0] reg_623__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_623(
    .clk(reg_623__clk),
    .in(reg_623__in),
    .out(reg_623__out)
  );

  //Wire declarations for instance 'reg_624' (Module coreir_reg)
  wire  reg_624__clk;
  wire [15:0] reg_624__in;
  wire [15:0] reg_624__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_624(
    .clk(reg_624__clk),
    .in(reg_624__in),
    .out(reg_624__out)
  );

  //Wire declarations for instance 'reg_625' (Module coreir_reg)
  wire  reg_625__clk;
  wire [15:0] reg_625__in;
  wire [15:0] reg_625__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_625(
    .clk(reg_625__clk),
    .in(reg_625__in),
    .out(reg_625__out)
  );

  //Wire declarations for instance 'reg_626' (Module coreir_reg)
  wire  reg_626__clk;
  wire [15:0] reg_626__in;
  wire [15:0] reg_626__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_626(
    .clk(reg_626__clk),
    .in(reg_626__in),
    .out(reg_626__out)
  );

  //Wire declarations for instance 'reg_627' (Module coreir_reg)
  wire  reg_627__clk;
  wire [15:0] reg_627__in;
  wire [15:0] reg_627__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_627(
    .clk(reg_627__clk),
    .in(reg_627__in),
    .out(reg_627__out)
  );

  //Wire declarations for instance 'reg_628' (Module coreir_reg)
  wire  reg_628__clk;
  wire [15:0] reg_628__in;
  wire [15:0] reg_628__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_628(
    .clk(reg_628__clk),
    .in(reg_628__in),
    .out(reg_628__out)
  );

  //Wire declarations for instance 'reg_629' (Module coreir_reg)
  wire  reg_629__clk;
  wire [15:0] reg_629__in;
  wire [15:0] reg_629__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_629(
    .clk(reg_629__clk),
    .in(reg_629__in),
    .out(reg_629__out)
  );

  //Wire declarations for instance 'reg_63' (Module coreir_reg)
  wire  reg_63__clk;
  wire [15:0] reg_63__in;
  wire [15:0] reg_63__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_63(
    .clk(reg_63__clk),
    .in(reg_63__in),
    .out(reg_63__out)
  );

  //Wire declarations for instance 'reg_630' (Module coreir_reg)
  wire  reg_630__clk;
  wire [15:0] reg_630__in;
  wire [15:0] reg_630__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_630(
    .clk(reg_630__clk),
    .in(reg_630__in),
    .out(reg_630__out)
  );

  //Wire declarations for instance 'reg_631' (Module coreir_reg)
  wire  reg_631__clk;
  wire [15:0] reg_631__in;
  wire [15:0] reg_631__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_631(
    .clk(reg_631__clk),
    .in(reg_631__in),
    .out(reg_631__out)
  );

  //Wire declarations for instance 'reg_632' (Module coreir_reg)
  wire  reg_632__clk;
  wire [15:0] reg_632__in;
  wire [15:0] reg_632__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_632(
    .clk(reg_632__clk),
    .in(reg_632__in),
    .out(reg_632__out)
  );

  //Wire declarations for instance 'reg_633' (Module coreir_reg)
  wire  reg_633__clk;
  wire [15:0] reg_633__in;
  wire [15:0] reg_633__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_633(
    .clk(reg_633__clk),
    .in(reg_633__in),
    .out(reg_633__out)
  );

  //Wire declarations for instance 'reg_634' (Module coreir_reg)
  wire  reg_634__clk;
  wire [15:0] reg_634__in;
  wire [15:0] reg_634__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_634(
    .clk(reg_634__clk),
    .in(reg_634__in),
    .out(reg_634__out)
  );

  //Wire declarations for instance 'reg_635' (Module coreir_reg)
  wire  reg_635__clk;
  wire [15:0] reg_635__in;
  wire [15:0] reg_635__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_635(
    .clk(reg_635__clk),
    .in(reg_635__in),
    .out(reg_635__out)
  );

  //Wire declarations for instance 'reg_636' (Module coreir_reg)
  wire  reg_636__clk;
  wire [15:0] reg_636__in;
  wire [15:0] reg_636__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_636(
    .clk(reg_636__clk),
    .in(reg_636__in),
    .out(reg_636__out)
  );

  //Wire declarations for instance 'reg_637' (Module coreir_reg)
  wire  reg_637__clk;
  wire [15:0] reg_637__in;
  wire [15:0] reg_637__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_637(
    .clk(reg_637__clk),
    .in(reg_637__in),
    .out(reg_637__out)
  );

  //Wire declarations for instance 'reg_638' (Module coreir_reg)
  wire  reg_638__clk;
  wire [15:0] reg_638__in;
  wire [15:0] reg_638__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_638(
    .clk(reg_638__clk),
    .in(reg_638__in),
    .out(reg_638__out)
  );

  //Wire declarations for instance 'reg_639' (Module coreir_reg)
  wire  reg_639__clk;
  wire [15:0] reg_639__in;
  wire [15:0] reg_639__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_639(
    .clk(reg_639__clk),
    .in(reg_639__in),
    .out(reg_639__out)
  );

  //Wire declarations for instance 'reg_64' (Module coreir_reg)
  wire  reg_64__clk;
  wire [15:0] reg_64__in;
  wire [15:0] reg_64__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_64(
    .clk(reg_64__clk),
    .in(reg_64__in),
    .out(reg_64__out)
  );

  //Wire declarations for instance 'reg_640' (Module coreir_reg)
  wire  reg_640__clk;
  wire [15:0] reg_640__in;
  wire [15:0] reg_640__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_640(
    .clk(reg_640__clk),
    .in(reg_640__in),
    .out(reg_640__out)
  );

  //Wire declarations for instance 'reg_641' (Module coreir_reg)
  wire  reg_641__clk;
  wire [15:0] reg_641__in;
  wire [15:0] reg_641__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_641(
    .clk(reg_641__clk),
    .in(reg_641__in),
    .out(reg_641__out)
  );

  //Wire declarations for instance 'reg_642' (Module coreir_reg)
  wire  reg_642__clk;
  wire [15:0] reg_642__in;
  wire [15:0] reg_642__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_642(
    .clk(reg_642__clk),
    .in(reg_642__in),
    .out(reg_642__out)
  );

  //Wire declarations for instance 'reg_643' (Module coreir_reg)
  wire  reg_643__clk;
  wire [15:0] reg_643__in;
  wire [15:0] reg_643__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_643(
    .clk(reg_643__clk),
    .in(reg_643__in),
    .out(reg_643__out)
  );

  //Wire declarations for instance 'reg_644' (Module coreir_reg)
  wire  reg_644__clk;
  wire [15:0] reg_644__in;
  wire [15:0] reg_644__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_644(
    .clk(reg_644__clk),
    .in(reg_644__in),
    .out(reg_644__out)
  );

  //Wire declarations for instance 'reg_645' (Module coreir_reg)
  wire  reg_645__clk;
  wire [15:0] reg_645__in;
  wire [15:0] reg_645__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_645(
    .clk(reg_645__clk),
    .in(reg_645__in),
    .out(reg_645__out)
  );

  //Wire declarations for instance 'reg_646' (Module coreir_reg)
  wire  reg_646__clk;
  wire [15:0] reg_646__in;
  wire [15:0] reg_646__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_646(
    .clk(reg_646__clk),
    .in(reg_646__in),
    .out(reg_646__out)
  );

  //Wire declarations for instance 'reg_647' (Module coreir_reg)
  wire  reg_647__clk;
  wire [15:0] reg_647__in;
  wire [15:0] reg_647__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_647(
    .clk(reg_647__clk),
    .in(reg_647__in),
    .out(reg_647__out)
  );

  //Wire declarations for instance 'reg_648' (Module coreir_reg)
  wire  reg_648__clk;
  wire [15:0] reg_648__in;
  wire [15:0] reg_648__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_648(
    .clk(reg_648__clk),
    .in(reg_648__in),
    .out(reg_648__out)
  );

  //Wire declarations for instance 'reg_649' (Module coreir_reg)
  wire  reg_649__clk;
  wire [15:0] reg_649__in;
  wire [15:0] reg_649__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_649(
    .clk(reg_649__clk),
    .in(reg_649__in),
    .out(reg_649__out)
  );

  //Wire declarations for instance 'reg_65' (Module coreir_reg)
  wire  reg_65__clk;
  wire [15:0] reg_65__in;
  wire [15:0] reg_65__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_65(
    .clk(reg_65__clk),
    .in(reg_65__in),
    .out(reg_65__out)
  );

  //Wire declarations for instance 'reg_650' (Module coreir_reg)
  wire  reg_650__clk;
  wire [15:0] reg_650__in;
  wire [15:0] reg_650__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_650(
    .clk(reg_650__clk),
    .in(reg_650__in),
    .out(reg_650__out)
  );

  //Wire declarations for instance 'reg_651' (Module coreir_reg)
  wire  reg_651__clk;
  wire [15:0] reg_651__in;
  wire [15:0] reg_651__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_651(
    .clk(reg_651__clk),
    .in(reg_651__in),
    .out(reg_651__out)
  );

  //Wire declarations for instance 'reg_652' (Module coreir_reg)
  wire  reg_652__clk;
  wire [15:0] reg_652__in;
  wire [15:0] reg_652__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_652(
    .clk(reg_652__clk),
    .in(reg_652__in),
    .out(reg_652__out)
  );

  //Wire declarations for instance 'reg_653' (Module coreir_reg)
  wire  reg_653__clk;
  wire [15:0] reg_653__in;
  wire [15:0] reg_653__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_653(
    .clk(reg_653__clk),
    .in(reg_653__in),
    .out(reg_653__out)
  );

  //Wire declarations for instance 'reg_654' (Module coreir_reg)
  wire  reg_654__clk;
  wire [15:0] reg_654__in;
  wire [15:0] reg_654__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_654(
    .clk(reg_654__clk),
    .in(reg_654__in),
    .out(reg_654__out)
  );

  //Wire declarations for instance 'reg_655' (Module coreir_reg)
  wire  reg_655__clk;
  wire [15:0] reg_655__in;
  wire [15:0] reg_655__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_655(
    .clk(reg_655__clk),
    .in(reg_655__in),
    .out(reg_655__out)
  );

  //Wire declarations for instance 'reg_656' (Module coreir_reg)
  wire  reg_656__clk;
  wire [15:0] reg_656__in;
  wire [15:0] reg_656__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_656(
    .clk(reg_656__clk),
    .in(reg_656__in),
    .out(reg_656__out)
  );

  //Wire declarations for instance 'reg_657' (Module coreir_reg)
  wire  reg_657__clk;
  wire [15:0] reg_657__in;
  wire [15:0] reg_657__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_657(
    .clk(reg_657__clk),
    .in(reg_657__in),
    .out(reg_657__out)
  );

  //Wire declarations for instance 'reg_658' (Module coreir_reg)
  wire  reg_658__clk;
  wire [15:0] reg_658__in;
  wire [15:0] reg_658__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_658(
    .clk(reg_658__clk),
    .in(reg_658__in),
    .out(reg_658__out)
  );

  //Wire declarations for instance 'reg_659' (Module coreir_reg)
  wire  reg_659__clk;
  wire [15:0] reg_659__in;
  wire [15:0] reg_659__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_659(
    .clk(reg_659__clk),
    .in(reg_659__in),
    .out(reg_659__out)
  );

  //Wire declarations for instance 'reg_66' (Module coreir_reg)
  wire  reg_66__clk;
  wire [15:0] reg_66__in;
  wire [15:0] reg_66__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_66(
    .clk(reg_66__clk),
    .in(reg_66__in),
    .out(reg_66__out)
  );

  //Wire declarations for instance 'reg_660' (Module coreir_reg)
  wire  reg_660__clk;
  wire [15:0] reg_660__in;
  wire [15:0] reg_660__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_660(
    .clk(reg_660__clk),
    .in(reg_660__in),
    .out(reg_660__out)
  );

  //Wire declarations for instance 'reg_661' (Module coreir_reg)
  wire  reg_661__clk;
  wire [15:0] reg_661__in;
  wire [15:0] reg_661__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_661(
    .clk(reg_661__clk),
    .in(reg_661__in),
    .out(reg_661__out)
  );

  //Wire declarations for instance 'reg_662' (Module coreir_reg)
  wire  reg_662__clk;
  wire [15:0] reg_662__in;
  wire [15:0] reg_662__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_662(
    .clk(reg_662__clk),
    .in(reg_662__in),
    .out(reg_662__out)
  );

  //Wire declarations for instance 'reg_663' (Module coreir_reg)
  wire  reg_663__clk;
  wire [15:0] reg_663__in;
  wire [15:0] reg_663__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_663(
    .clk(reg_663__clk),
    .in(reg_663__in),
    .out(reg_663__out)
  );

  //Wire declarations for instance 'reg_664' (Module coreir_reg)
  wire  reg_664__clk;
  wire [15:0] reg_664__in;
  wire [15:0] reg_664__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_664(
    .clk(reg_664__clk),
    .in(reg_664__in),
    .out(reg_664__out)
  );

  //Wire declarations for instance 'reg_665' (Module coreir_reg)
  wire  reg_665__clk;
  wire [15:0] reg_665__in;
  wire [15:0] reg_665__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_665(
    .clk(reg_665__clk),
    .in(reg_665__in),
    .out(reg_665__out)
  );

  //Wire declarations for instance 'reg_666' (Module coreir_reg)
  wire  reg_666__clk;
  wire [15:0] reg_666__in;
  wire [15:0] reg_666__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_666(
    .clk(reg_666__clk),
    .in(reg_666__in),
    .out(reg_666__out)
  );

  //Wire declarations for instance 'reg_667' (Module coreir_reg)
  wire  reg_667__clk;
  wire [15:0] reg_667__in;
  wire [15:0] reg_667__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_667(
    .clk(reg_667__clk),
    .in(reg_667__in),
    .out(reg_667__out)
  );

  //Wire declarations for instance 'reg_668' (Module coreir_reg)
  wire  reg_668__clk;
  wire [15:0] reg_668__in;
  wire [15:0] reg_668__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_668(
    .clk(reg_668__clk),
    .in(reg_668__in),
    .out(reg_668__out)
  );

  //Wire declarations for instance 'reg_669' (Module coreir_reg)
  wire  reg_669__clk;
  wire [15:0] reg_669__in;
  wire [15:0] reg_669__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_669(
    .clk(reg_669__clk),
    .in(reg_669__in),
    .out(reg_669__out)
  );

  //Wire declarations for instance 'reg_67' (Module coreir_reg)
  wire  reg_67__clk;
  wire [15:0] reg_67__in;
  wire [15:0] reg_67__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_67(
    .clk(reg_67__clk),
    .in(reg_67__in),
    .out(reg_67__out)
  );

  //Wire declarations for instance 'reg_670' (Module coreir_reg)
  wire  reg_670__clk;
  wire [15:0] reg_670__in;
  wire [15:0] reg_670__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_670(
    .clk(reg_670__clk),
    .in(reg_670__in),
    .out(reg_670__out)
  );

  //Wire declarations for instance 'reg_671' (Module coreir_reg)
  wire  reg_671__clk;
  wire [15:0] reg_671__in;
  wire [15:0] reg_671__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_671(
    .clk(reg_671__clk),
    .in(reg_671__in),
    .out(reg_671__out)
  );

  //Wire declarations for instance 'reg_672' (Module coreir_reg)
  wire  reg_672__clk;
  wire [15:0] reg_672__in;
  wire [15:0] reg_672__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_672(
    .clk(reg_672__clk),
    .in(reg_672__in),
    .out(reg_672__out)
  );

  //Wire declarations for instance 'reg_673' (Module coreir_reg)
  wire  reg_673__clk;
  wire [15:0] reg_673__in;
  wire [15:0] reg_673__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_673(
    .clk(reg_673__clk),
    .in(reg_673__in),
    .out(reg_673__out)
  );

  //Wire declarations for instance 'reg_674' (Module coreir_reg)
  wire  reg_674__clk;
  wire [15:0] reg_674__in;
  wire [15:0] reg_674__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_674(
    .clk(reg_674__clk),
    .in(reg_674__in),
    .out(reg_674__out)
  );

  //Wire declarations for instance 'reg_675' (Module coreir_reg)
  wire  reg_675__clk;
  wire [15:0] reg_675__in;
  wire [15:0] reg_675__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_675(
    .clk(reg_675__clk),
    .in(reg_675__in),
    .out(reg_675__out)
  );

  //Wire declarations for instance 'reg_676' (Module coreir_reg)
  wire  reg_676__clk;
  wire [15:0] reg_676__in;
  wire [15:0] reg_676__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_676(
    .clk(reg_676__clk),
    .in(reg_676__in),
    .out(reg_676__out)
  );

  //Wire declarations for instance 'reg_677' (Module coreir_reg)
  wire  reg_677__clk;
  wire [15:0] reg_677__in;
  wire [15:0] reg_677__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_677(
    .clk(reg_677__clk),
    .in(reg_677__in),
    .out(reg_677__out)
  );

  //Wire declarations for instance 'reg_678' (Module coreir_reg)
  wire  reg_678__clk;
  wire [15:0] reg_678__in;
  wire [15:0] reg_678__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_678(
    .clk(reg_678__clk),
    .in(reg_678__in),
    .out(reg_678__out)
  );

  //Wire declarations for instance 'reg_679' (Module coreir_reg)
  wire  reg_679__clk;
  wire [15:0] reg_679__in;
  wire [15:0] reg_679__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_679(
    .clk(reg_679__clk),
    .in(reg_679__in),
    .out(reg_679__out)
  );

  //Wire declarations for instance 'reg_68' (Module coreir_reg)
  wire  reg_68__clk;
  wire [15:0] reg_68__in;
  wire [15:0] reg_68__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_68(
    .clk(reg_68__clk),
    .in(reg_68__in),
    .out(reg_68__out)
  );

  //Wire declarations for instance 'reg_680' (Module coreir_reg)
  wire  reg_680__clk;
  wire [15:0] reg_680__in;
  wire [15:0] reg_680__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_680(
    .clk(reg_680__clk),
    .in(reg_680__in),
    .out(reg_680__out)
  );

  //Wire declarations for instance 'reg_681' (Module coreir_reg)
  wire  reg_681__clk;
  wire [15:0] reg_681__in;
  wire [15:0] reg_681__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_681(
    .clk(reg_681__clk),
    .in(reg_681__in),
    .out(reg_681__out)
  );

  //Wire declarations for instance 'reg_682' (Module coreir_reg)
  wire  reg_682__clk;
  wire [15:0] reg_682__in;
  wire [15:0] reg_682__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_682(
    .clk(reg_682__clk),
    .in(reg_682__in),
    .out(reg_682__out)
  );

  //Wire declarations for instance 'reg_683' (Module coreir_reg)
  wire  reg_683__clk;
  wire [15:0] reg_683__in;
  wire [15:0] reg_683__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_683(
    .clk(reg_683__clk),
    .in(reg_683__in),
    .out(reg_683__out)
  );

  //Wire declarations for instance 'reg_684' (Module coreir_reg)
  wire  reg_684__clk;
  wire [15:0] reg_684__in;
  wire [15:0] reg_684__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_684(
    .clk(reg_684__clk),
    .in(reg_684__in),
    .out(reg_684__out)
  );

  //Wire declarations for instance 'reg_685' (Module coreir_reg)
  wire  reg_685__clk;
  wire [15:0] reg_685__in;
  wire [15:0] reg_685__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_685(
    .clk(reg_685__clk),
    .in(reg_685__in),
    .out(reg_685__out)
  );

  //Wire declarations for instance 'reg_686' (Module coreir_reg)
  wire  reg_686__clk;
  wire [15:0] reg_686__in;
  wire [15:0] reg_686__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_686(
    .clk(reg_686__clk),
    .in(reg_686__in),
    .out(reg_686__out)
  );

  //Wire declarations for instance 'reg_687' (Module coreir_reg)
  wire  reg_687__clk;
  wire [15:0] reg_687__in;
  wire [15:0] reg_687__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_687(
    .clk(reg_687__clk),
    .in(reg_687__in),
    .out(reg_687__out)
  );

  //Wire declarations for instance 'reg_688' (Module coreir_reg)
  wire  reg_688__clk;
  wire [15:0] reg_688__in;
  wire [15:0] reg_688__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_688(
    .clk(reg_688__clk),
    .in(reg_688__in),
    .out(reg_688__out)
  );

  //Wire declarations for instance 'reg_689' (Module coreir_reg)
  wire  reg_689__clk;
  wire [15:0] reg_689__in;
  wire [15:0] reg_689__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_689(
    .clk(reg_689__clk),
    .in(reg_689__in),
    .out(reg_689__out)
  );

  //Wire declarations for instance 'reg_69' (Module coreir_reg)
  wire  reg_69__clk;
  wire [15:0] reg_69__in;
  wire [15:0] reg_69__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_69(
    .clk(reg_69__clk),
    .in(reg_69__in),
    .out(reg_69__out)
  );

  //Wire declarations for instance 'reg_690' (Module coreir_reg)
  wire  reg_690__clk;
  wire [15:0] reg_690__in;
  wire [15:0] reg_690__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_690(
    .clk(reg_690__clk),
    .in(reg_690__in),
    .out(reg_690__out)
  );

  //Wire declarations for instance 'reg_691' (Module coreir_reg)
  wire  reg_691__clk;
  wire [15:0] reg_691__in;
  wire [15:0] reg_691__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_691(
    .clk(reg_691__clk),
    .in(reg_691__in),
    .out(reg_691__out)
  );

  //Wire declarations for instance 'reg_692' (Module coreir_reg)
  wire  reg_692__clk;
  wire [15:0] reg_692__in;
  wire [15:0] reg_692__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_692(
    .clk(reg_692__clk),
    .in(reg_692__in),
    .out(reg_692__out)
  );

  //Wire declarations for instance 'reg_693' (Module coreir_reg)
  wire  reg_693__clk;
  wire [15:0] reg_693__in;
  wire [15:0] reg_693__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_693(
    .clk(reg_693__clk),
    .in(reg_693__in),
    .out(reg_693__out)
  );

  //Wire declarations for instance 'reg_694' (Module coreir_reg)
  wire  reg_694__clk;
  wire [15:0] reg_694__in;
  wire [15:0] reg_694__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_694(
    .clk(reg_694__clk),
    .in(reg_694__in),
    .out(reg_694__out)
  );

  //Wire declarations for instance 'reg_695' (Module coreir_reg)
  wire  reg_695__clk;
  wire [15:0] reg_695__in;
  wire [15:0] reg_695__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_695(
    .clk(reg_695__clk),
    .in(reg_695__in),
    .out(reg_695__out)
  );

  //Wire declarations for instance 'reg_696' (Module coreir_reg)
  wire  reg_696__clk;
  wire [15:0] reg_696__in;
  wire [15:0] reg_696__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_696(
    .clk(reg_696__clk),
    .in(reg_696__in),
    .out(reg_696__out)
  );

  //Wire declarations for instance 'reg_697' (Module coreir_reg)
  wire  reg_697__clk;
  wire [15:0] reg_697__in;
  wire [15:0] reg_697__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_697(
    .clk(reg_697__clk),
    .in(reg_697__in),
    .out(reg_697__out)
  );

  //Wire declarations for instance 'reg_698' (Module coreir_reg)
  wire  reg_698__clk;
  wire [15:0] reg_698__in;
  wire [15:0] reg_698__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_698(
    .clk(reg_698__clk),
    .in(reg_698__in),
    .out(reg_698__out)
  );

  //Wire declarations for instance 'reg_699' (Module coreir_reg)
  wire  reg_699__clk;
  wire [15:0] reg_699__in;
  wire [15:0] reg_699__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_699(
    .clk(reg_699__clk),
    .in(reg_699__in),
    .out(reg_699__out)
  );

  //Wire declarations for instance 'reg_7' (Module coreir_reg)
  wire  reg_7__clk;
  wire [15:0] reg_7__in;
  wire [15:0] reg_7__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_7(
    .clk(reg_7__clk),
    .in(reg_7__in),
    .out(reg_7__out)
  );

  //Wire declarations for instance 'reg_70' (Module coreir_reg)
  wire  reg_70__clk;
  wire [15:0] reg_70__in;
  wire [15:0] reg_70__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_70(
    .clk(reg_70__clk),
    .in(reg_70__in),
    .out(reg_70__out)
  );

  //Wire declarations for instance 'reg_700' (Module coreir_reg)
  wire  reg_700__clk;
  wire [15:0] reg_700__in;
  wire [15:0] reg_700__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_700(
    .clk(reg_700__clk),
    .in(reg_700__in),
    .out(reg_700__out)
  );

  //Wire declarations for instance 'reg_701' (Module coreir_reg)
  wire  reg_701__clk;
  wire [15:0] reg_701__in;
  wire [15:0] reg_701__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_701(
    .clk(reg_701__clk),
    .in(reg_701__in),
    .out(reg_701__out)
  );

  //Wire declarations for instance 'reg_702' (Module coreir_reg)
  wire  reg_702__clk;
  wire [15:0] reg_702__in;
  wire [15:0] reg_702__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_702(
    .clk(reg_702__clk),
    .in(reg_702__in),
    .out(reg_702__out)
  );

  //Wire declarations for instance 'reg_703' (Module coreir_reg)
  wire  reg_703__clk;
  wire [15:0] reg_703__in;
  wire [15:0] reg_703__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_703(
    .clk(reg_703__clk),
    .in(reg_703__in),
    .out(reg_703__out)
  );

  //Wire declarations for instance 'reg_704' (Module coreir_reg)
  wire  reg_704__clk;
  wire [15:0] reg_704__in;
  wire [15:0] reg_704__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_704(
    .clk(reg_704__clk),
    .in(reg_704__in),
    .out(reg_704__out)
  );

  //Wire declarations for instance 'reg_705' (Module coreir_reg)
  wire  reg_705__clk;
  wire [15:0] reg_705__in;
  wire [15:0] reg_705__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_705(
    .clk(reg_705__clk),
    .in(reg_705__in),
    .out(reg_705__out)
  );

  //Wire declarations for instance 'reg_706' (Module coreir_reg)
  wire  reg_706__clk;
  wire [15:0] reg_706__in;
  wire [15:0] reg_706__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_706(
    .clk(reg_706__clk),
    .in(reg_706__in),
    .out(reg_706__out)
  );

  //Wire declarations for instance 'reg_707' (Module coreir_reg)
  wire  reg_707__clk;
  wire [15:0] reg_707__in;
  wire [15:0] reg_707__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_707(
    .clk(reg_707__clk),
    .in(reg_707__in),
    .out(reg_707__out)
  );

  //Wire declarations for instance 'reg_708' (Module coreir_reg)
  wire  reg_708__clk;
  wire [15:0] reg_708__in;
  wire [15:0] reg_708__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_708(
    .clk(reg_708__clk),
    .in(reg_708__in),
    .out(reg_708__out)
  );

  //Wire declarations for instance 'reg_709' (Module coreir_reg)
  wire  reg_709__clk;
  wire [15:0] reg_709__in;
  wire [15:0] reg_709__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_709(
    .clk(reg_709__clk),
    .in(reg_709__in),
    .out(reg_709__out)
  );

  //Wire declarations for instance 'reg_71' (Module coreir_reg)
  wire  reg_71__clk;
  wire [15:0] reg_71__in;
  wire [15:0] reg_71__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_71(
    .clk(reg_71__clk),
    .in(reg_71__in),
    .out(reg_71__out)
  );

  //Wire declarations for instance 'reg_710' (Module coreir_reg)
  wire  reg_710__clk;
  wire [15:0] reg_710__in;
  wire [15:0] reg_710__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_710(
    .clk(reg_710__clk),
    .in(reg_710__in),
    .out(reg_710__out)
  );

  //Wire declarations for instance 'reg_711' (Module coreir_reg)
  wire  reg_711__clk;
  wire [15:0] reg_711__in;
  wire [15:0] reg_711__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_711(
    .clk(reg_711__clk),
    .in(reg_711__in),
    .out(reg_711__out)
  );

  //Wire declarations for instance 'reg_712' (Module coreir_reg)
  wire  reg_712__clk;
  wire [15:0] reg_712__in;
  wire [15:0] reg_712__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_712(
    .clk(reg_712__clk),
    .in(reg_712__in),
    .out(reg_712__out)
  );

  //Wire declarations for instance 'reg_713' (Module coreir_reg)
  wire  reg_713__clk;
  wire [15:0] reg_713__in;
  wire [15:0] reg_713__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_713(
    .clk(reg_713__clk),
    .in(reg_713__in),
    .out(reg_713__out)
  );

  //Wire declarations for instance 'reg_714' (Module coreir_reg)
  wire  reg_714__clk;
  wire [15:0] reg_714__in;
  wire [15:0] reg_714__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_714(
    .clk(reg_714__clk),
    .in(reg_714__in),
    .out(reg_714__out)
  );

  //Wire declarations for instance 'reg_715' (Module coreir_reg)
  wire  reg_715__clk;
  wire [15:0] reg_715__in;
  wire [15:0] reg_715__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_715(
    .clk(reg_715__clk),
    .in(reg_715__in),
    .out(reg_715__out)
  );

  //Wire declarations for instance 'reg_716' (Module coreir_reg)
  wire  reg_716__clk;
  wire [15:0] reg_716__in;
  wire [15:0] reg_716__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_716(
    .clk(reg_716__clk),
    .in(reg_716__in),
    .out(reg_716__out)
  );

  //Wire declarations for instance 'reg_717' (Module coreir_reg)
  wire  reg_717__clk;
  wire [15:0] reg_717__in;
  wire [15:0] reg_717__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_717(
    .clk(reg_717__clk),
    .in(reg_717__in),
    .out(reg_717__out)
  );

  //Wire declarations for instance 'reg_718' (Module coreir_reg)
  wire  reg_718__clk;
  wire [15:0] reg_718__in;
  wire [15:0] reg_718__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_718(
    .clk(reg_718__clk),
    .in(reg_718__in),
    .out(reg_718__out)
  );

  //Wire declarations for instance 'reg_719' (Module coreir_reg)
  wire  reg_719__clk;
  wire [15:0] reg_719__in;
  wire [15:0] reg_719__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_719(
    .clk(reg_719__clk),
    .in(reg_719__in),
    .out(reg_719__out)
  );

  //Wire declarations for instance 'reg_72' (Module coreir_reg)
  wire  reg_72__clk;
  wire [15:0] reg_72__in;
  wire [15:0] reg_72__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_72(
    .clk(reg_72__clk),
    .in(reg_72__in),
    .out(reg_72__out)
  );

  //Wire declarations for instance 'reg_720' (Module coreir_reg)
  wire  reg_720__clk;
  wire [15:0] reg_720__in;
  wire [15:0] reg_720__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_720(
    .clk(reg_720__clk),
    .in(reg_720__in),
    .out(reg_720__out)
  );

  //Wire declarations for instance 'reg_721' (Module coreir_reg)
  wire  reg_721__clk;
  wire [15:0] reg_721__in;
  wire [15:0] reg_721__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_721(
    .clk(reg_721__clk),
    .in(reg_721__in),
    .out(reg_721__out)
  );

  //Wire declarations for instance 'reg_722' (Module coreir_reg)
  wire  reg_722__clk;
  wire [15:0] reg_722__in;
  wire [15:0] reg_722__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_722(
    .clk(reg_722__clk),
    .in(reg_722__in),
    .out(reg_722__out)
  );

  //Wire declarations for instance 'reg_723' (Module coreir_reg)
  wire  reg_723__clk;
  wire [15:0] reg_723__in;
  wire [15:0] reg_723__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_723(
    .clk(reg_723__clk),
    .in(reg_723__in),
    .out(reg_723__out)
  );

  //Wire declarations for instance 'reg_724' (Module coreir_reg)
  wire  reg_724__clk;
  wire [15:0] reg_724__in;
  wire [15:0] reg_724__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_724(
    .clk(reg_724__clk),
    .in(reg_724__in),
    .out(reg_724__out)
  );

  //Wire declarations for instance 'reg_725' (Module coreir_reg)
  wire  reg_725__clk;
  wire [15:0] reg_725__in;
  wire [15:0] reg_725__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_725(
    .clk(reg_725__clk),
    .in(reg_725__in),
    .out(reg_725__out)
  );

  //Wire declarations for instance 'reg_726' (Module coreir_reg)
  wire  reg_726__clk;
  wire [15:0] reg_726__in;
  wire [15:0] reg_726__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_726(
    .clk(reg_726__clk),
    .in(reg_726__in),
    .out(reg_726__out)
  );

  //Wire declarations for instance 'reg_727' (Module coreir_reg)
  wire  reg_727__clk;
  wire [15:0] reg_727__in;
  wire [15:0] reg_727__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_727(
    .clk(reg_727__clk),
    .in(reg_727__in),
    .out(reg_727__out)
  );

  //Wire declarations for instance 'reg_728' (Module coreir_reg)
  wire  reg_728__clk;
  wire [15:0] reg_728__in;
  wire [15:0] reg_728__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_728(
    .clk(reg_728__clk),
    .in(reg_728__in),
    .out(reg_728__out)
  );

  //Wire declarations for instance 'reg_729' (Module coreir_reg)
  wire  reg_729__clk;
  wire [15:0] reg_729__in;
  wire [15:0] reg_729__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_729(
    .clk(reg_729__clk),
    .in(reg_729__in),
    .out(reg_729__out)
  );

  //Wire declarations for instance 'reg_73' (Module coreir_reg)
  wire  reg_73__clk;
  wire [15:0] reg_73__in;
  wire [15:0] reg_73__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_73(
    .clk(reg_73__clk),
    .in(reg_73__in),
    .out(reg_73__out)
  );

  //Wire declarations for instance 'reg_730' (Module coreir_reg)
  wire  reg_730__clk;
  wire [15:0] reg_730__in;
  wire [15:0] reg_730__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_730(
    .clk(reg_730__clk),
    .in(reg_730__in),
    .out(reg_730__out)
  );

  //Wire declarations for instance 'reg_731' (Module coreir_reg)
  wire  reg_731__clk;
  wire [15:0] reg_731__in;
  wire [15:0] reg_731__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_731(
    .clk(reg_731__clk),
    .in(reg_731__in),
    .out(reg_731__out)
  );

  //Wire declarations for instance 'reg_732' (Module coreir_reg)
  wire  reg_732__clk;
  wire [15:0] reg_732__in;
  wire [15:0] reg_732__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_732(
    .clk(reg_732__clk),
    .in(reg_732__in),
    .out(reg_732__out)
  );

  //Wire declarations for instance 'reg_733' (Module coreir_reg)
  wire  reg_733__clk;
  wire [15:0] reg_733__in;
  wire [15:0] reg_733__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_733(
    .clk(reg_733__clk),
    .in(reg_733__in),
    .out(reg_733__out)
  );

  //Wire declarations for instance 'reg_734' (Module coreir_reg)
  wire  reg_734__clk;
  wire [15:0] reg_734__in;
  wire [15:0] reg_734__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_734(
    .clk(reg_734__clk),
    .in(reg_734__in),
    .out(reg_734__out)
  );

  //Wire declarations for instance 'reg_735' (Module coreir_reg)
  wire  reg_735__clk;
  wire [15:0] reg_735__in;
  wire [15:0] reg_735__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_735(
    .clk(reg_735__clk),
    .in(reg_735__in),
    .out(reg_735__out)
  );

  //Wire declarations for instance 'reg_736' (Module coreir_reg)
  wire  reg_736__clk;
  wire [15:0] reg_736__in;
  wire [15:0] reg_736__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_736(
    .clk(reg_736__clk),
    .in(reg_736__in),
    .out(reg_736__out)
  );

  //Wire declarations for instance 'reg_737' (Module coreir_reg)
  wire  reg_737__clk;
  wire [15:0] reg_737__in;
  wire [15:0] reg_737__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_737(
    .clk(reg_737__clk),
    .in(reg_737__in),
    .out(reg_737__out)
  );

  //Wire declarations for instance 'reg_738' (Module coreir_reg)
  wire  reg_738__clk;
  wire [15:0] reg_738__in;
  wire [15:0] reg_738__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_738(
    .clk(reg_738__clk),
    .in(reg_738__in),
    .out(reg_738__out)
  );

  //Wire declarations for instance 'reg_739' (Module coreir_reg)
  wire  reg_739__clk;
  wire [15:0] reg_739__in;
  wire [15:0] reg_739__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_739(
    .clk(reg_739__clk),
    .in(reg_739__in),
    .out(reg_739__out)
  );

  //Wire declarations for instance 'reg_74' (Module coreir_reg)
  wire  reg_74__clk;
  wire [15:0] reg_74__in;
  wire [15:0] reg_74__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_74(
    .clk(reg_74__clk),
    .in(reg_74__in),
    .out(reg_74__out)
  );

  //Wire declarations for instance 'reg_740' (Module coreir_reg)
  wire  reg_740__clk;
  wire [15:0] reg_740__in;
  wire [15:0] reg_740__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_740(
    .clk(reg_740__clk),
    .in(reg_740__in),
    .out(reg_740__out)
  );

  //Wire declarations for instance 'reg_741' (Module coreir_reg)
  wire  reg_741__clk;
  wire [15:0] reg_741__in;
  wire [15:0] reg_741__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_741(
    .clk(reg_741__clk),
    .in(reg_741__in),
    .out(reg_741__out)
  );

  //Wire declarations for instance 'reg_742' (Module coreir_reg)
  wire  reg_742__clk;
  wire [15:0] reg_742__in;
  wire [15:0] reg_742__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_742(
    .clk(reg_742__clk),
    .in(reg_742__in),
    .out(reg_742__out)
  );

  //Wire declarations for instance 'reg_743' (Module coreir_reg)
  wire  reg_743__clk;
  wire [15:0] reg_743__in;
  wire [15:0] reg_743__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_743(
    .clk(reg_743__clk),
    .in(reg_743__in),
    .out(reg_743__out)
  );

  //Wire declarations for instance 'reg_744' (Module coreir_reg)
  wire  reg_744__clk;
  wire [15:0] reg_744__in;
  wire [15:0] reg_744__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_744(
    .clk(reg_744__clk),
    .in(reg_744__in),
    .out(reg_744__out)
  );

  //Wire declarations for instance 'reg_745' (Module coreir_reg)
  wire  reg_745__clk;
  wire [15:0] reg_745__in;
  wire [15:0] reg_745__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_745(
    .clk(reg_745__clk),
    .in(reg_745__in),
    .out(reg_745__out)
  );

  //Wire declarations for instance 'reg_746' (Module coreir_reg)
  wire  reg_746__clk;
  wire [15:0] reg_746__in;
  wire [15:0] reg_746__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_746(
    .clk(reg_746__clk),
    .in(reg_746__in),
    .out(reg_746__out)
  );

  //Wire declarations for instance 'reg_747' (Module coreir_reg)
  wire  reg_747__clk;
  wire [15:0] reg_747__in;
  wire [15:0] reg_747__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_747(
    .clk(reg_747__clk),
    .in(reg_747__in),
    .out(reg_747__out)
  );

  //Wire declarations for instance 'reg_748' (Module coreir_reg)
  wire  reg_748__clk;
  wire [15:0] reg_748__in;
  wire [15:0] reg_748__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_748(
    .clk(reg_748__clk),
    .in(reg_748__in),
    .out(reg_748__out)
  );

  //Wire declarations for instance 'reg_749' (Module coreir_reg)
  wire  reg_749__clk;
  wire [15:0] reg_749__in;
  wire [15:0] reg_749__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_749(
    .clk(reg_749__clk),
    .in(reg_749__in),
    .out(reg_749__out)
  );

  //Wire declarations for instance 'reg_75' (Module coreir_reg)
  wire  reg_75__clk;
  wire [15:0] reg_75__in;
  wire [15:0] reg_75__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_75(
    .clk(reg_75__clk),
    .in(reg_75__in),
    .out(reg_75__out)
  );

  //Wire declarations for instance 'reg_750' (Module coreir_reg)
  wire  reg_750__clk;
  wire [15:0] reg_750__in;
  wire [15:0] reg_750__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_750(
    .clk(reg_750__clk),
    .in(reg_750__in),
    .out(reg_750__out)
  );

  //Wire declarations for instance 'reg_751' (Module coreir_reg)
  wire  reg_751__clk;
  wire [15:0] reg_751__in;
  wire [15:0] reg_751__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_751(
    .clk(reg_751__clk),
    .in(reg_751__in),
    .out(reg_751__out)
  );

  //Wire declarations for instance 'reg_752' (Module coreir_reg)
  wire  reg_752__clk;
  wire [15:0] reg_752__in;
  wire [15:0] reg_752__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_752(
    .clk(reg_752__clk),
    .in(reg_752__in),
    .out(reg_752__out)
  );

  //Wire declarations for instance 'reg_753' (Module coreir_reg)
  wire  reg_753__clk;
  wire [15:0] reg_753__in;
  wire [15:0] reg_753__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_753(
    .clk(reg_753__clk),
    .in(reg_753__in),
    .out(reg_753__out)
  );

  //Wire declarations for instance 'reg_754' (Module coreir_reg)
  wire  reg_754__clk;
  wire [15:0] reg_754__in;
  wire [15:0] reg_754__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_754(
    .clk(reg_754__clk),
    .in(reg_754__in),
    .out(reg_754__out)
  );

  //Wire declarations for instance 'reg_755' (Module coreir_reg)
  wire  reg_755__clk;
  wire [15:0] reg_755__in;
  wire [15:0] reg_755__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_755(
    .clk(reg_755__clk),
    .in(reg_755__in),
    .out(reg_755__out)
  );

  //Wire declarations for instance 'reg_756' (Module coreir_reg)
  wire  reg_756__clk;
  wire [15:0] reg_756__in;
  wire [15:0] reg_756__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_756(
    .clk(reg_756__clk),
    .in(reg_756__in),
    .out(reg_756__out)
  );

  //Wire declarations for instance 'reg_757' (Module coreir_reg)
  wire  reg_757__clk;
  wire [15:0] reg_757__in;
  wire [15:0] reg_757__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_757(
    .clk(reg_757__clk),
    .in(reg_757__in),
    .out(reg_757__out)
  );

  //Wire declarations for instance 'reg_758' (Module coreir_reg)
  wire  reg_758__clk;
  wire [15:0] reg_758__in;
  wire [15:0] reg_758__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_758(
    .clk(reg_758__clk),
    .in(reg_758__in),
    .out(reg_758__out)
  );

  //Wire declarations for instance 'reg_759' (Module coreir_reg)
  wire  reg_759__clk;
  wire [15:0] reg_759__in;
  wire [15:0] reg_759__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_759(
    .clk(reg_759__clk),
    .in(reg_759__in),
    .out(reg_759__out)
  );

  //Wire declarations for instance 'reg_76' (Module coreir_reg)
  wire  reg_76__clk;
  wire [15:0] reg_76__in;
  wire [15:0] reg_76__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_76(
    .clk(reg_76__clk),
    .in(reg_76__in),
    .out(reg_76__out)
  );

  //Wire declarations for instance 'reg_760' (Module coreir_reg)
  wire  reg_760__clk;
  wire [15:0] reg_760__in;
  wire [15:0] reg_760__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_760(
    .clk(reg_760__clk),
    .in(reg_760__in),
    .out(reg_760__out)
  );

  //Wire declarations for instance 'reg_761' (Module coreir_reg)
  wire  reg_761__clk;
  wire [15:0] reg_761__in;
  wire [15:0] reg_761__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_761(
    .clk(reg_761__clk),
    .in(reg_761__in),
    .out(reg_761__out)
  );

  //Wire declarations for instance 'reg_762' (Module coreir_reg)
  wire  reg_762__clk;
  wire [15:0] reg_762__in;
  wire [15:0] reg_762__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_762(
    .clk(reg_762__clk),
    .in(reg_762__in),
    .out(reg_762__out)
  );

  //Wire declarations for instance 'reg_763' (Module coreir_reg)
  wire  reg_763__clk;
  wire [15:0] reg_763__in;
  wire [15:0] reg_763__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_763(
    .clk(reg_763__clk),
    .in(reg_763__in),
    .out(reg_763__out)
  );

  //Wire declarations for instance 'reg_764' (Module coreir_reg)
  wire  reg_764__clk;
  wire [15:0] reg_764__in;
  wire [15:0] reg_764__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_764(
    .clk(reg_764__clk),
    .in(reg_764__in),
    .out(reg_764__out)
  );

  //Wire declarations for instance 'reg_765' (Module coreir_reg)
  wire  reg_765__clk;
  wire [15:0] reg_765__in;
  wire [15:0] reg_765__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_765(
    .clk(reg_765__clk),
    .in(reg_765__in),
    .out(reg_765__out)
  );

  //Wire declarations for instance 'reg_766' (Module coreir_reg)
  wire  reg_766__clk;
  wire [15:0] reg_766__in;
  wire [15:0] reg_766__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_766(
    .clk(reg_766__clk),
    .in(reg_766__in),
    .out(reg_766__out)
  );

  //Wire declarations for instance 'reg_767' (Module coreir_reg)
  wire  reg_767__clk;
  wire [15:0] reg_767__in;
  wire [15:0] reg_767__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_767(
    .clk(reg_767__clk),
    .in(reg_767__in),
    .out(reg_767__out)
  );

  //Wire declarations for instance 'reg_768' (Module coreir_reg)
  wire  reg_768__clk;
  wire [15:0] reg_768__in;
  wire [15:0] reg_768__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_768(
    .clk(reg_768__clk),
    .in(reg_768__in),
    .out(reg_768__out)
  );

  //Wire declarations for instance 'reg_769' (Module coreir_reg)
  wire  reg_769__clk;
  wire [15:0] reg_769__in;
  wire [15:0] reg_769__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_769(
    .clk(reg_769__clk),
    .in(reg_769__in),
    .out(reg_769__out)
  );

  //Wire declarations for instance 'reg_77' (Module coreir_reg)
  wire  reg_77__clk;
  wire [15:0] reg_77__in;
  wire [15:0] reg_77__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_77(
    .clk(reg_77__clk),
    .in(reg_77__in),
    .out(reg_77__out)
  );

  //Wire declarations for instance 'reg_770' (Module coreir_reg)
  wire  reg_770__clk;
  wire [15:0] reg_770__in;
  wire [15:0] reg_770__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_770(
    .clk(reg_770__clk),
    .in(reg_770__in),
    .out(reg_770__out)
  );

  //Wire declarations for instance 'reg_771' (Module coreir_reg)
  wire  reg_771__clk;
  wire [15:0] reg_771__in;
  wire [15:0] reg_771__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_771(
    .clk(reg_771__clk),
    .in(reg_771__in),
    .out(reg_771__out)
  );

  //Wire declarations for instance 'reg_772' (Module coreir_reg)
  wire  reg_772__clk;
  wire [15:0] reg_772__in;
  wire [15:0] reg_772__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_772(
    .clk(reg_772__clk),
    .in(reg_772__in),
    .out(reg_772__out)
  );

  //Wire declarations for instance 'reg_773' (Module coreir_reg)
  wire  reg_773__clk;
  wire [15:0] reg_773__in;
  wire [15:0] reg_773__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_773(
    .clk(reg_773__clk),
    .in(reg_773__in),
    .out(reg_773__out)
  );

  //Wire declarations for instance 'reg_774' (Module coreir_reg)
  wire  reg_774__clk;
  wire [15:0] reg_774__in;
  wire [15:0] reg_774__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_774(
    .clk(reg_774__clk),
    .in(reg_774__in),
    .out(reg_774__out)
  );

  //Wire declarations for instance 'reg_775' (Module coreir_reg)
  wire  reg_775__clk;
  wire [15:0] reg_775__in;
  wire [15:0] reg_775__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_775(
    .clk(reg_775__clk),
    .in(reg_775__in),
    .out(reg_775__out)
  );

  //Wire declarations for instance 'reg_776' (Module coreir_reg)
  wire  reg_776__clk;
  wire [15:0] reg_776__in;
  wire [15:0] reg_776__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_776(
    .clk(reg_776__clk),
    .in(reg_776__in),
    .out(reg_776__out)
  );

  //Wire declarations for instance 'reg_777' (Module coreir_reg)
  wire  reg_777__clk;
  wire [15:0] reg_777__in;
  wire [15:0] reg_777__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_777(
    .clk(reg_777__clk),
    .in(reg_777__in),
    .out(reg_777__out)
  );

  //Wire declarations for instance 'reg_778' (Module coreir_reg)
  wire  reg_778__clk;
  wire [15:0] reg_778__in;
  wire [15:0] reg_778__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_778(
    .clk(reg_778__clk),
    .in(reg_778__in),
    .out(reg_778__out)
  );

  //Wire declarations for instance 'reg_779' (Module coreir_reg)
  wire  reg_779__clk;
  wire [15:0] reg_779__in;
  wire [15:0] reg_779__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_779(
    .clk(reg_779__clk),
    .in(reg_779__in),
    .out(reg_779__out)
  );

  //Wire declarations for instance 'reg_78' (Module coreir_reg)
  wire  reg_78__clk;
  wire [15:0] reg_78__in;
  wire [15:0] reg_78__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_78(
    .clk(reg_78__clk),
    .in(reg_78__in),
    .out(reg_78__out)
  );

  //Wire declarations for instance 'reg_780' (Module coreir_reg)
  wire  reg_780__clk;
  wire [15:0] reg_780__in;
  wire [15:0] reg_780__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_780(
    .clk(reg_780__clk),
    .in(reg_780__in),
    .out(reg_780__out)
  );

  //Wire declarations for instance 'reg_781' (Module coreir_reg)
  wire  reg_781__clk;
  wire [15:0] reg_781__in;
  wire [15:0] reg_781__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_781(
    .clk(reg_781__clk),
    .in(reg_781__in),
    .out(reg_781__out)
  );

  //Wire declarations for instance 'reg_782' (Module coreir_reg)
  wire  reg_782__clk;
  wire [15:0] reg_782__in;
  wire [15:0] reg_782__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_782(
    .clk(reg_782__clk),
    .in(reg_782__in),
    .out(reg_782__out)
  );

  //Wire declarations for instance 'reg_783' (Module coreir_reg)
  wire  reg_783__clk;
  wire [15:0] reg_783__in;
  wire [15:0] reg_783__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_783(
    .clk(reg_783__clk),
    .in(reg_783__in),
    .out(reg_783__out)
  );

  //Wire declarations for instance 'reg_784' (Module coreir_reg)
  wire  reg_784__clk;
  wire [15:0] reg_784__in;
  wire [15:0] reg_784__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_784(
    .clk(reg_784__clk),
    .in(reg_784__in),
    .out(reg_784__out)
  );

  //Wire declarations for instance 'reg_785' (Module coreir_reg)
  wire  reg_785__clk;
  wire [15:0] reg_785__in;
  wire [15:0] reg_785__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_785(
    .clk(reg_785__clk),
    .in(reg_785__in),
    .out(reg_785__out)
  );

  //Wire declarations for instance 'reg_786' (Module coreir_reg)
  wire  reg_786__clk;
  wire [15:0] reg_786__in;
  wire [15:0] reg_786__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_786(
    .clk(reg_786__clk),
    .in(reg_786__in),
    .out(reg_786__out)
  );

  //Wire declarations for instance 'reg_787' (Module coreir_reg)
  wire  reg_787__clk;
  wire [15:0] reg_787__in;
  wire [15:0] reg_787__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_787(
    .clk(reg_787__clk),
    .in(reg_787__in),
    .out(reg_787__out)
  );

  //Wire declarations for instance 'reg_788' (Module coreir_reg)
  wire  reg_788__clk;
  wire [15:0] reg_788__in;
  wire [15:0] reg_788__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_788(
    .clk(reg_788__clk),
    .in(reg_788__in),
    .out(reg_788__out)
  );

  //Wire declarations for instance 'reg_789' (Module coreir_reg)
  wire  reg_789__clk;
  wire [15:0] reg_789__in;
  wire [15:0] reg_789__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_789(
    .clk(reg_789__clk),
    .in(reg_789__in),
    .out(reg_789__out)
  );

  //Wire declarations for instance 'reg_79' (Module coreir_reg)
  wire  reg_79__clk;
  wire [15:0] reg_79__in;
  wire [15:0] reg_79__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_79(
    .clk(reg_79__clk),
    .in(reg_79__in),
    .out(reg_79__out)
  );

  //Wire declarations for instance 'reg_790' (Module coreir_reg)
  wire  reg_790__clk;
  wire [15:0] reg_790__in;
  wire [15:0] reg_790__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_790(
    .clk(reg_790__clk),
    .in(reg_790__in),
    .out(reg_790__out)
  );

  //Wire declarations for instance 'reg_791' (Module coreir_reg)
  wire  reg_791__clk;
  wire [15:0] reg_791__in;
  wire [15:0] reg_791__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_791(
    .clk(reg_791__clk),
    .in(reg_791__in),
    .out(reg_791__out)
  );

  //Wire declarations for instance 'reg_792' (Module coreir_reg)
  wire  reg_792__clk;
  wire [15:0] reg_792__in;
  wire [15:0] reg_792__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_792(
    .clk(reg_792__clk),
    .in(reg_792__in),
    .out(reg_792__out)
  );

  //Wire declarations for instance 'reg_793' (Module coreir_reg)
  wire  reg_793__clk;
  wire [15:0] reg_793__in;
  wire [15:0] reg_793__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_793(
    .clk(reg_793__clk),
    .in(reg_793__in),
    .out(reg_793__out)
  );

  //Wire declarations for instance 'reg_794' (Module coreir_reg)
  wire  reg_794__clk;
  wire [15:0] reg_794__in;
  wire [15:0] reg_794__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_794(
    .clk(reg_794__clk),
    .in(reg_794__in),
    .out(reg_794__out)
  );

  //Wire declarations for instance 'reg_795' (Module coreir_reg)
  wire  reg_795__clk;
  wire [15:0] reg_795__in;
  wire [15:0] reg_795__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_795(
    .clk(reg_795__clk),
    .in(reg_795__in),
    .out(reg_795__out)
  );

  //Wire declarations for instance 'reg_796' (Module coreir_reg)
  wire  reg_796__clk;
  wire [15:0] reg_796__in;
  wire [15:0] reg_796__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_796(
    .clk(reg_796__clk),
    .in(reg_796__in),
    .out(reg_796__out)
  );

  //Wire declarations for instance 'reg_797' (Module coreir_reg)
  wire  reg_797__clk;
  wire [15:0] reg_797__in;
  wire [15:0] reg_797__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_797(
    .clk(reg_797__clk),
    .in(reg_797__in),
    .out(reg_797__out)
  );

  //Wire declarations for instance 'reg_798' (Module coreir_reg)
  wire  reg_798__clk;
  wire [15:0] reg_798__in;
  wire [15:0] reg_798__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_798(
    .clk(reg_798__clk),
    .in(reg_798__in),
    .out(reg_798__out)
  );

  //Wire declarations for instance 'reg_799' (Module coreir_reg)
  wire  reg_799__clk;
  wire [15:0] reg_799__in;
  wire [15:0] reg_799__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_799(
    .clk(reg_799__clk),
    .in(reg_799__in),
    .out(reg_799__out)
  );

  //Wire declarations for instance 'reg_8' (Module coreir_reg)
  wire  reg_8__clk;
  wire [15:0] reg_8__in;
  wire [15:0] reg_8__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_8(
    .clk(reg_8__clk),
    .in(reg_8__in),
    .out(reg_8__out)
  );

  //Wire declarations for instance 'reg_80' (Module coreir_reg)
  wire  reg_80__clk;
  wire [15:0] reg_80__in;
  wire [15:0] reg_80__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_80(
    .clk(reg_80__clk),
    .in(reg_80__in),
    .out(reg_80__out)
  );

  //Wire declarations for instance 'reg_800' (Module coreir_reg)
  wire  reg_800__clk;
  wire [15:0] reg_800__in;
  wire [15:0] reg_800__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_800(
    .clk(reg_800__clk),
    .in(reg_800__in),
    .out(reg_800__out)
  );

  //Wire declarations for instance 'reg_801' (Module coreir_reg)
  wire  reg_801__clk;
  wire [15:0] reg_801__in;
  wire [15:0] reg_801__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_801(
    .clk(reg_801__clk),
    .in(reg_801__in),
    .out(reg_801__out)
  );

  //Wire declarations for instance 'reg_802' (Module coreir_reg)
  wire  reg_802__clk;
  wire [15:0] reg_802__in;
  wire [15:0] reg_802__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_802(
    .clk(reg_802__clk),
    .in(reg_802__in),
    .out(reg_802__out)
  );

  //Wire declarations for instance 'reg_803' (Module coreir_reg)
  wire  reg_803__clk;
  wire [15:0] reg_803__in;
  wire [15:0] reg_803__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_803(
    .clk(reg_803__clk),
    .in(reg_803__in),
    .out(reg_803__out)
  );

  //Wire declarations for instance 'reg_804' (Module coreir_reg)
  wire  reg_804__clk;
  wire [15:0] reg_804__in;
  wire [15:0] reg_804__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_804(
    .clk(reg_804__clk),
    .in(reg_804__in),
    .out(reg_804__out)
  );

  //Wire declarations for instance 'reg_805' (Module coreir_reg)
  wire  reg_805__clk;
  wire [15:0] reg_805__in;
  wire [15:0] reg_805__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_805(
    .clk(reg_805__clk),
    .in(reg_805__in),
    .out(reg_805__out)
  );

  //Wire declarations for instance 'reg_806' (Module coreir_reg)
  wire  reg_806__clk;
  wire [15:0] reg_806__in;
  wire [15:0] reg_806__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_806(
    .clk(reg_806__clk),
    .in(reg_806__in),
    .out(reg_806__out)
  );

  //Wire declarations for instance 'reg_807' (Module coreir_reg)
  wire  reg_807__clk;
  wire [15:0] reg_807__in;
  wire [15:0] reg_807__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_807(
    .clk(reg_807__clk),
    .in(reg_807__in),
    .out(reg_807__out)
  );

  //Wire declarations for instance 'reg_808' (Module coreir_reg)
  wire  reg_808__clk;
  wire [15:0] reg_808__in;
  wire [15:0] reg_808__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_808(
    .clk(reg_808__clk),
    .in(reg_808__in),
    .out(reg_808__out)
  );

  //Wire declarations for instance 'reg_809' (Module coreir_reg)
  wire  reg_809__clk;
  wire [15:0] reg_809__in;
  wire [15:0] reg_809__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_809(
    .clk(reg_809__clk),
    .in(reg_809__in),
    .out(reg_809__out)
  );

  //Wire declarations for instance 'reg_81' (Module coreir_reg)
  wire  reg_81__clk;
  wire [15:0] reg_81__in;
  wire [15:0] reg_81__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_81(
    .clk(reg_81__clk),
    .in(reg_81__in),
    .out(reg_81__out)
  );

  //Wire declarations for instance 'reg_810' (Module coreir_reg)
  wire  reg_810__clk;
  wire [15:0] reg_810__in;
  wire [15:0] reg_810__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_810(
    .clk(reg_810__clk),
    .in(reg_810__in),
    .out(reg_810__out)
  );

  //Wire declarations for instance 'reg_811' (Module coreir_reg)
  wire  reg_811__clk;
  wire [15:0] reg_811__in;
  wire [15:0] reg_811__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_811(
    .clk(reg_811__clk),
    .in(reg_811__in),
    .out(reg_811__out)
  );

  //Wire declarations for instance 'reg_812' (Module coreir_reg)
  wire  reg_812__clk;
  wire [15:0] reg_812__in;
  wire [15:0] reg_812__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_812(
    .clk(reg_812__clk),
    .in(reg_812__in),
    .out(reg_812__out)
  );

  //Wire declarations for instance 'reg_813' (Module coreir_reg)
  wire  reg_813__clk;
  wire [15:0] reg_813__in;
  wire [15:0] reg_813__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_813(
    .clk(reg_813__clk),
    .in(reg_813__in),
    .out(reg_813__out)
  );

  //Wire declarations for instance 'reg_814' (Module coreir_reg)
  wire  reg_814__clk;
  wire [15:0] reg_814__in;
  wire [15:0] reg_814__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_814(
    .clk(reg_814__clk),
    .in(reg_814__in),
    .out(reg_814__out)
  );

  //Wire declarations for instance 'reg_815' (Module coreir_reg)
  wire  reg_815__clk;
  wire [15:0] reg_815__in;
  wire [15:0] reg_815__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_815(
    .clk(reg_815__clk),
    .in(reg_815__in),
    .out(reg_815__out)
  );

  //Wire declarations for instance 'reg_816' (Module coreir_reg)
  wire  reg_816__clk;
  wire [15:0] reg_816__in;
  wire [15:0] reg_816__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_816(
    .clk(reg_816__clk),
    .in(reg_816__in),
    .out(reg_816__out)
  );

  //Wire declarations for instance 'reg_817' (Module coreir_reg)
  wire  reg_817__clk;
  wire [15:0] reg_817__in;
  wire [15:0] reg_817__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_817(
    .clk(reg_817__clk),
    .in(reg_817__in),
    .out(reg_817__out)
  );

  //Wire declarations for instance 'reg_818' (Module coreir_reg)
  wire  reg_818__clk;
  wire [15:0] reg_818__in;
  wire [15:0] reg_818__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_818(
    .clk(reg_818__clk),
    .in(reg_818__in),
    .out(reg_818__out)
  );

  //Wire declarations for instance 'reg_819' (Module coreir_reg)
  wire  reg_819__clk;
  wire [15:0] reg_819__in;
  wire [15:0] reg_819__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_819(
    .clk(reg_819__clk),
    .in(reg_819__in),
    .out(reg_819__out)
  );

  //Wire declarations for instance 'reg_82' (Module coreir_reg)
  wire  reg_82__clk;
  wire [15:0] reg_82__in;
  wire [15:0] reg_82__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_82(
    .clk(reg_82__clk),
    .in(reg_82__in),
    .out(reg_82__out)
  );

  //Wire declarations for instance 'reg_820' (Module coreir_reg)
  wire  reg_820__clk;
  wire [15:0] reg_820__in;
  wire [15:0] reg_820__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_820(
    .clk(reg_820__clk),
    .in(reg_820__in),
    .out(reg_820__out)
  );

  //Wire declarations for instance 'reg_821' (Module coreir_reg)
  wire  reg_821__clk;
  wire [15:0] reg_821__in;
  wire [15:0] reg_821__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_821(
    .clk(reg_821__clk),
    .in(reg_821__in),
    .out(reg_821__out)
  );

  //Wire declarations for instance 'reg_822' (Module coreir_reg)
  wire  reg_822__clk;
  wire [15:0] reg_822__in;
  wire [15:0] reg_822__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_822(
    .clk(reg_822__clk),
    .in(reg_822__in),
    .out(reg_822__out)
  );

  //Wire declarations for instance 'reg_823' (Module coreir_reg)
  wire  reg_823__clk;
  wire [15:0] reg_823__in;
  wire [15:0] reg_823__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_823(
    .clk(reg_823__clk),
    .in(reg_823__in),
    .out(reg_823__out)
  );

  //Wire declarations for instance 'reg_824' (Module coreir_reg)
  wire  reg_824__clk;
  wire [15:0] reg_824__in;
  wire [15:0] reg_824__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_824(
    .clk(reg_824__clk),
    .in(reg_824__in),
    .out(reg_824__out)
  );

  //Wire declarations for instance 'reg_825' (Module coreir_reg)
  wire  reg_825__clk;
  wire [15:0] reg_825__in;
  wire [15:0] reg_825__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_825(
    .clk(reg_825__clk),
    .in(reg_825__in),
    .out(reg_825__out)
  );

  //Wire declarations for instance 'reg_826' (Module coreir_reg)
  wire  reg_826__clk;
  wire [15:0] reg_826__in;
  wire [15:0] reg_826__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_826(
    .clk(reg_826__clk),
    .in(reg_826__in),
    .out(reg_826__out)
  );

  //Wire declarations for instance 'reg_827' (Module coreir_reg)
  wire  reg_827__clk;
  wire [15:0] reg_827__in;
  wire [15:0] reg_827__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_827(
    .clk(reg_827__clk),
    .in(reg_827__in),
    .out(reg_827__out)
  );

  //Wire declarations for instance 'reg_828' (Module coreir_reg)
  wire  reg_828__clk;
  wire [15:0] reg_828__in;
  wire [15:0] reg_828__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_828(
    .clk(reg_828__clk),
    .in(reg_828__in),
    .out(reg_828__out)
  );

  //Wire declarations for instance 'reg_829' (Module coreir_reg)
  wire  reg_829__clk;
  wire [15:0] reg_829__in;
  wire [15:0] reg_829__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_829(
    .clk(reg_829__clk),
    .in(reg_829__in),
    .out(reg_829__out)
  );

  //Wire declarations for instance 'reg_83' (Module coreir_reg)
  wire  reg_83__clk;
  wire [15:0] reg_83__in;
  wire [15:0] reg_83__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_83(
    .clk(reg_83__clk),
    .in(reg_83__in),
    .out(reg_83__out)
  );

  //Wire declarations for instance 'reg_830' (Module coreir_reg)
  wire  reg_830__clk;
  wire [15:0] reg_830__in;
  wire [15:0] reg_830__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_830(
    .clk(reg_830__clk),
    .in(reg_830__in),
    .out(reg_830__out)
  );

  //Wire declarations for instance 'reg_831' (Module coreir_reg)
  wire  reg_831__clk;
  wire [15:0] reg_831__in;
  wire [15:0] reg_831__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_831(
    .clk(reg_831__clk),
    .in(reg_831__in),
    .out(reg_831__out)
  );

  //Wire declarations for instance 'reg_832' (Module coreir_reg)
  wire  reg_832__clk;
  wire [15:0] reg_832__in;
  wire [15:0] reg_832__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_832(
    .clk(reg_832__clk),
    .in(reg_832__in),
    .out(reg_832__out)
  );

  //Wire declarations for instance 'reg_833' (Module coreir_reg)
  wire  reg_833__clk;
  wire [15:0] reg_833__in;
  wire [15:0] reg_833__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_833(
    .clk(reg_833__clk),
    .in(reg_833__in),
    .out(reg_833__out)
  );

  //Wire declarations for instance 'reg_834' (Module coreir_reg)
  wire  reg_834__clk;
  wire [15:0] reg_834__in;
  wire [15:0] reg_834__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_834(
    .clk(reg_834__clk),
    .in(reg_834__in),
    .out(reg_834__out)
  );

  //Wire declarations for instance 'reg_835' (Module coreir_reg)
  wire  reg_835__clk;
  wire [15:0] reg_835__in;
  wire [15:0] reg_835__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_835(
    .clk(reg_835__clk),
    .in(reg_835__in),
    .out(reg_835__out)
  );

  //Wire declarations for instance 'reg_836' (Module coreir_reg)
  wire  reg_836__clk;
  wire [15:0] reg_836__in;
  wire [15:0] reg_836__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_836(
    .clk(reg_836__clk),
    .in(reg_836__in),
    .out(reg_836__out)
  );

  //Wire declarations for instance 'reg_837' (Module coreir_reg)
  wire  reg_837__clk;
  wire [15:0] reg_837__in;
  wire [15:0] reg_837__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_837(
    .clk(reg_837__clk),
    .in(reg_837__in),
    .out(reg_837__out)
  );

  //Wire declarations for instance 'reg_838' (Module coreir_reg)
  wire  reg_838__clk;
  wire [15:0] reg_838__in;
  wire [15:0] reg_838__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_838(
    .clk(reg_838__clk),
    .in(reg_838__in),
    .out(reg_838__out)
  );

  //Wire declarations for instance 'reg_839' (Module coreir_reg)
  wire  reg_839__clk;
  wire [15:0] reg_839__in;
  wire [15:0] reg_839__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_839(
    .clk(reg_839__clk),
    .in(reg_839__in),
    .out(reg_839__out)
  );

  //Wire declarations for instance 'reg_84' (Module coreir_reg)
  wire  reg_84__clk;
  wire [15:0] reg_84__in;
  wire [15:0] reg_84__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_84(
    .clk(reg_84__clk),
    .in(reg_84__in),
    .out(reg_84__out)
  );

  //Wire declarations for instance 'reg_840' (Module coreir_reg)
  wire  reg_840__clk;
  wire [15:0] reg_840__in;
  wire [15:0] reg_840__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_840(
    .clk(reg_840__clk),
    .in(reg_840__in),
    .out(reg_840__out)
  );

  //Wire declarations for instance 'reg_841' (Module coreir_reg)
  wire  reg_841__clk;
  wire [15:0] reg_841__in;
  wire [15:0] reg_841__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_841(
    .clk(reg_841__clk),
    .in(reg_841__in),
    .out(reg_841__out)
  );

  //Wire declarations for instance 'reg_842' (Module coreir_reg)
  wire  reg_842__clk;
  wire [15:0] reg_842__in;
  wire [15:0] reg_842__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_842(
    .clk(reg_842__clk),
    .in(reg_842__in),
    .out(reg_842__out)
  );

  //Wire declarations for instance 'reg_843' (Module coreir_reg)
  wire  reg_843__clk;
  wire [15:0] reg_843__in;
  wire [15:0] reg_843__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_843(
    .clk(reg_843__clk),
    .in(reg_843__in),
    .out(reg_843__out)
  );

  //Wire declarations for instance 'reg_844' (Module coreir_reg)
  wire  reg_844__clk;
  wire [15:0] reg_844__in;
  wire [15:0] reg_844__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_844(
    .clk(reg_844__clk),
    .in(reg_844__in),
    .out(reg_844__out)
  );

  //Wire declarations for instance 'reg_845' (Module coreir_reg)
  wire  reg_845__clk;
  wire [15:0] reg_845__in;
  wire [15:0] reg_845__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_845(
    .clk(reg_845__clk),
    .in(reg_845__in),
    .out(reg_845__out)
  );

  //Wire declarations for instance 'reg_846' (Module coreir_reg)
  wire  reg_846__clk;
  wire [15:0] reg_846__in;
  wire [15:0] reg_846__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_846(
    .clk(reg_846__clk),
    .in(reg_846__in),
    .out(reg_846__out)
  );

  //Wire declarations for instance 'reg_847' (Module coreir_reg)
  wire  reg_847__clk;
  wire [15:0] reg_847__in;
  wire [15:0] reg_847__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_847(
    .clk(reg_847__clk),
    .in(reg_847__in),
    .out(reg_847__out)
  );

  //Wire declarations for instance 'reg_848' (Module coreir_reg)
  wire  reg_848__clk;
  wire [15:0] reg_848__in;
  wire [15:0] reg_848__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_848(
    .clk(reg_848__clk),
    .in(reg_848__in),
    .out(reg_848__out)
  );

  //Wire declarations for instance 'reg_849' (Module coreir_reg)
  wire  reg_849__clk;
  wire [15:0] reg_849__in;
  wire [15:0] reg_849__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_849(
    .clk(reg_849__clk),
    .in(reg_849__in),
    .out(reg_849__out)
  );

  //Wire declarations for instance 'reg_85' (Module coreir_reg)
  wire  reg_85__clk;
  wire [15:0] reg_85__in;
  wire [15:0] reg_85__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_85(
    .clk(reg_85__clk),
    .in(reg_85__in),
    .out(reg_85__out)
  );

  //Wire declarations for instance 'reg_850' (Module coreir_reg)
  wire  reg_850__clk;
  wire [15:0] reg_850__in;
  wire [15:0] reg_850__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_850(
    .clk(reg_850__clk),
    .in(reg_850__in),
    .out(reg_850__out)
  );

  //Wire declarations for instance 'reg_851' (Module coreir_reg)
  wire  reg_851__clk;
  wire [15:0] reg_851__in;
  wire [15:0] reg_851__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_851(
    .clk(reg_851__clk),
    .in(reg_851__in),
    .out(reg_851__out)
  );

  //Wire declarations for instance 'reg_852' (Module coreir_reg)
  wire  reg_852__clk;
  wire [15:0] reg_852__in;
  wire [15:0] reg_852__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_852(
    .clk(reg_852__clk),
    .in(reg_852__in),
    .out(reg_852__out)
  );

  //Wire declarations for instance 'reg_853' (Module coreir_reg)
  wire  reg_853__clk;
  wire [15:0] reg_853__in;
  wire [15:0] reg_853__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_853(
    .clk(reg_853__clk),
    .in(reg_853__in),
    .out(reg_853__out)
  );

  //Wire declarations for instance 'reg_854' (Module coreir_reg)
  wire  reg_854__clk;
  wire [15:0] reg_854__in;
  wire [15:0] reg_854__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_854(
    .clk(reg_854__clk),
    .in(reg_854__in),
    .out(reg_854__out)
  );

  //Wire declarations for instance 'reg_855' (Module coreir_reg)
  wire  reg_855__clk;
  wire [15:0] reg_855__in;
  wire [15:0] reg_855__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_855(
    .clk(reg_855__clk),
    .in(reg_855__in),
    .out(reg_855__out)
  );

  //Wire declarations for instance 'reg_856' (Module coreir_reg)
  wire  reg_856__clk;
  wire [15:0] reg_856__in;
  wire [15:0] reg_856__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_856(
    .clk(reg_856__clk),
    .in(reg_856__in),
    .out(reg_856__out)
  );

  //Wire declarations for instance 'reg_857' (Module coreir_reg)
  wire  reg_857__clk;
  wire [15:0] reg_857__in;
  wire [15:0] reg_857__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_857(
    .clk(reg_857__clk),
    .in(reg_857__in),
    .out(reg_857__out)
  );

  //Wire declarations for instance 'reg_858' (Module coreir_reg)
  wire  reg_858__clk;
  wire [15:0] reg_858__in;
  wire [15:0] reg_858__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_858(
    .clk(reg_858__clk),
    .in(reg_858__in),
    .out(reg_858__out)
  );

  //Wire declarations for instance 'reg_859' (Module coreir_reg)
  wire  reg_859__clk;
  wire [15:0] reg_859__in;
  wire [15:0] reg_859__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_859(
    .clk(reg_859__clk),
    .in(reg_859__in),
    .out(reg_859__out)
  );

  //Wire declarations for instance 'reg_86' (Module coreir_reg)
  wire  reg_86__clk;
  wire [15:0] reg_86__in;
  wire [15:0] reg_86__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_86(
    .clk(reg_86__clk),
    .in(reg_86__in),
    .out(reg_86__out)
  );

  //Wire declarations for instance 'reg_860' (Module coreir_reg)
  wire  reg_860__clk;
  wire [15:0] reg_860__in;
  wire [15:0] reg_860__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_860(
    .clk(reg_860__clk),
    .in(reg_860__in),
    .out(reg_860__out)
  );

  //Wire declarations for instance 'reg_861' (Module coreir_reg)
  wire  reg_861__clk;
  wire [15:0] reg_861__in;
  wire [15:0] reg_861__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_861(
    .clk(reg_861__clk),
    .in(reg_861__in),
    .out(reg_861__out)
  );

  //Wire declarations for instance 'reg_862' (Module coreir_reg)
  wire  reg_862__clk;
  wire [15:0] reg_862__in;
  wire [15:0] reg_862__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_862(
    .clk(reg_862__clk),
    .in(reg_862__in),
    .out(reg_862__out)
  );

  //Wire declarations for instance 'reg_863' (Module coreir_reg)
  wire  reg_863__clk;
  wire [15:0] reg_863__in;
  wire [15:0] reg_863__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_863(
    .clk(reg_863__clk),
    .in(reg_863__in),
    .out(reg_863__out)
  );

  //Wire declarations for instance 'reg_864' (Module coreir_reg)
  wire  reg_864__clk;
  wire [15:0] reg_864__in;
  wire [15:0] reg_864__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_864(
    .clk(reg_864__clk),
    .in(reg_864__in),
    .out(reg_864__out)
  );

  //Wire declarations for instance 'reg_865' (Module coreir_reg)
  wire  reg_865__clk;
  wire [15:0] reg_865__in;
  wire [15:0] reg_865__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_865(
    .clk(reg_865__clk),
    .in(reg_865__in),
    .out(reg_865__out)
  );

  //Wire declarations for instance 'reg_866' (Module coreir_reg)
  wire  reg_866__clk;
  wire [15:0] reg_866__in;
  wire [15:0] reg_866__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_866(
    .clk(reg_866__clk),
    .in(reg_866__in),
    .out(reg_866__out)
  );

  //Wire declarations for instance 'reg_867' (Module coreir_reg)
  wire  reg_867__clk;
  wire [15:0] reg_867__in;
  wire [15:0] reg_867__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_867(
    .clk(reg_867__clk),
    .in(reg_867__in),
    .out(reg_867__out)
  );

  //Wire declarations for instance 'reg_868' (Module coreir_reg)
  wire  reg_868__clk;
  wire [15:0] reg_868__in;
  wire [15:0] reg_868__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_868(
    .clk(reg_868__clk),
    .in(reg_868__in),
    .out(reg_868__out)
  );

  //Wire declarations for instance 'reg_869' (Module coreir_reg)
  wire  reg_869__clk;
  wire [15:0] reg_869__in;
  wire [15:0] reg_869__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_869(
    .clk(reg_869__clk),
    .in(reg_869__in),
    .out(reg_869__out)
  );

  //Wire declarations for instance 'reg_87' (Module coreir_reg)
  wire  reg_87__clk;
  wire [15:0] reg_87__in;
  wire [15:0] reg_87__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_87(
    .clk(reg_87__clk),
    .in(reg_87__in),
    .out(reg_87__out)
  );

  //Wire declarations for instance 'reg_870' (Module coreir_reg)
  wire  reg_870__clk;
  wire [15:0] reg_870__in;
  wire [15:0] reg_870__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_870(
    .clk(reg_870__clk),
    .in(reg_870__in),
    .out(reg_870__out)
  );

  //Wire declarations for instance 'reg_871' (Module coreir_reg)
  wire  reg_871__clk;
  wire [15:0] reg_871__in;
  wire [15:0] reg_871__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_871(
    .clk(reg_871__clk),
    .in(reg_871__in),
    .out(reg_871__out)
  );

  //Wire declarations for instance 'reg_872' (Module coreir_reg)
  wire  reg_872__clk;
  wire [15:0] reg_872__in;
  wire [15:0] reg_872__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_872(
    .clk(reg_872__clk),
    .in(reg_872__in),
    .out(reg_872__out)
  );

  //Wire declarations for instance 'reg_873' (Module coreir_reg)
  wire  reg_873__clk;
  wire [15:0] reg_873__in;
  wire [15:0] reg_873__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_873(
    .clk(reg_873__clk),
    .in(reg_873__in),
    .out(reg_873__out)
  );

  //Wire declarations for instance 'reg_874' (Module coreir_reg)
  wire  reg_874__clk;
  wire [15:0] reg_874__in;
  wire [15:0] reg_874__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_874(
    .clk(reg_874__clk),
    .in(reg_874__in),
    .out(reg_874__out)
  );

  //Wire declarations for instance 'reg_875' (Module coreir_reg)
  wire  reg_875__clk;
  wire [15:0] reg_875__in;
  wire [15:0] reg_875__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_875(
    .clk(reg_875__clk),
    .in(reg_875__in),
    .out(reg_875__out)
  );

  //Wire declarations for instance 'reg_876' (Module coreir_reg)
  wire  reg_876__clk;
  wire [15:0] reg_876__in;
  wire [15:0] reg_876__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_876(
    .clk(reg_876__clk),
    .in(reg_876__in),
    .out(reg_876__out)
  );

  //Wire declarations for instance 'reg_877' (Module coreir_reg)
  wire  reg_877__clk;
  wire [15:0] reg_877__in;
  wire [15:0] reg_877__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_877(
    .clk(reg_877__clk),
    .in(reg_877__in),
    .out(reg_877__out)
  );

  //Wire declarations for instance 'reg_878' (Module coreir_reg)
  wire  reg_878__clk;
  wire [15:0] reg_878__in;
  wire [15:0] reg_878__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_878(
    .clk(reg_878__clk),
    .in(reg_878__in),
    .out(reg_878__out)
  );

  //Wire declarations for instance 'reg_879' (Module coreir_reg)
  wire  reg_879__clk;
  wire [15:0] reg_879__in;
  wire [15:0] reg_879__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_879(
    .clk(reg_879__clk),
    .in(reg_879__in),
    .out(reg_879__out)
  );

  //Wire declarations for instance 'reg_88' (Module coreir_reg)
  wire  reg_88__clk;
  wire [15:0] reg_88__in;
  wire [15:0] reg_88__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_88(
    .clk(reg_88__clk),
    .in(reg_88__in),
    .out(reg_88__out)
  );

  //Wire declarations for instance 'reg_880' (Module coreir_reg)
  wire  reg_880__clk;
  wire [15:0] reg_880__in;
  wire [15:0] reg_880__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_880(
    .clk(reg_880__clk),
    .in(reg_880__in),
    .out(reg_880__out)
  );

  //Wire declarations for instance 'reg_881' (Module coreir_reg)
  wire  reg_881__clk;
  wire [15:0] reg_881__in;
  wire [15:0] reg_881__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_881(
    .clk(reg_881__clk),
    .in(reg_881__in),
    .out(reg_881__out)
  );

  //Wire declarations for instance 'reg_882' (Module coreir_reg)
  wire  reg_882__clk;
  wire [15:0] reg_882__in;
  wire [15:0] reg_882__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_882(
    .clk(reg_882__clk),
    .in(reg_882__in),
    .out(reg_882__out)
  );

  //Wire declarations for instance 'reg_883' (Module coreir_reg)
  wire  reg_883__clk;
  wire [15:0] reg_883__in;
  wire [15:0] reg_883__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_883(
    .clk(reg_883__clk),
    .in(reg_883__in),
    .out(reg_883__out)
  );

  //Wire declarations for instance 'reg_884' (Module coreir_reg)
  wire  reg_884__clk;
  wire [15:0] reg_884__in;
  wire [15:0] reg_884__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_884(
    .clk(reg_884__clk),
    .in(reg_884__in),
    .out(reg_884__out)
  );

  //Wire declarations for instance 'reg_885' (Module coreir_reg)
  wire  reg_885__clk;
  wire [15:0] reg_885__in;
  wire [15:0] reg_885__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_885(
    .clk(reg_885__clk),
    .in(reg_885__in),
    .out(reg_885__out)
  );

  //Wire declarations for instance 'reg_886' (Module coreir_reg)
  wire  reg_886__clk;
  wire [15:0] reg_886__in;
  wire [15:0] reg_886__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_886(
    .clk(reg_886__clk),
    .in(reg_886__in),
    .out(reg_886__out)
  );

  //Wire declarations for instance 'reg_887' (Module coreir_reg)
  wire  reg_887__clk;
  wire [15:0] reg_887__in;
  wire [15:0] reg_887__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_887(
    .clk(reg_887__clk),
    .in(reg_887__in),
    .out(reg_887__out)
  );

  //Wire declarations for instance 'reg_888' (Module coreir_reg)
  wire  reg_888__clk;
  wire [15:0] reg_888__in;
  wire [15:0] reg_888__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_888(
    .clk(reg_888__clk),
    .in(reg_888__in),
    .out(reg_888__out)
  );

  //Wire declarations for instance 'reg_889' (Module coreir_reg)
  wire  reg_889__clk;
  wire [15:0] reg_889__in;
  wire [15:0] reg_889__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_889(
    .clk(reg_889__clk),
    .in(reg_889__in),
    .out(reg_889__out)
  );

  //Wire declarations for instance 'reg_89' (Module coreir_reg)
  wire  reg_89__clk;
  wire [15:0] reg_89__in;
  wire [15:0] reg_89__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_89(
    .clk(reg_89__clk),
    .in(reg_89__in),
    .out(reg_89__out)
  );

  //Wire declarations for instance 'reg_890' (Module coreir_reg)
  wire  reg_890__clk;
  wire [15:0] reg_890__in;
  wire [15:0] reg_890__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_890(
    .clk(reg_890__clk),
    .in(reg_890__in),
    .out(reg_890__out)
  );

  //Wire declarations for instance 'reg_891' (Module coreir_reg)
  wire  reg_891__clk;
  wire [15:0] reg_891__in;
  wire [15:0] reg_891__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_891(
    .clk(reg_891__clk),
    .in(reg_891__in),
    .out(reg_891__out)
  );

  //Wire declarations for instance 'reg_892' (Module coreir_reg)
  wire  reg_892__clk;
  wire [15:0] reg_892__in;
  wire [15:0] reg_892__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_892(
    .clk(reg_892__clk),
    .in(reg_892__in),
    .out(reg_892__out)
  );

  //Wire declarations for instance 'reg_893' (Module coreir_reg)
  wire  reg_893__clk;
  wire [15:0] reg_893__in;
  wire [15:0] reg_893__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_893(
    .clk(reg_893__clk),
    .in(reg_893__in),
    .out(reg_893__out)
  );

  //Wire declarations for instance 'reg_894' (Module coreir_reg)
  wire  reg_894__clk;
  wire [15:0] reg_894__in;
  wire [15:0] reg_894__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_894(
    .clk(reg_894__clk),
    .in(reg_894__in),
    .out(reg_894__out)
  );

  //Wire declarations for instance 'reg_895' (Module coreir_reg)
  wire  reg_895__clk;
  wire [15:0] reg_895__in;
  wire [15:0] reg_895__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_895(
    .clk(reg_895__clk),
    .in(reg_895__in),
    .out(reg_895__out)
  );

  //Wire declarations for instance 'reg_896' (Module coreir_reg)
  wire  reg_896__clk;
  wire [15:0] reg_896__in;
  wire [15:0] reg_896__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_896(
    .clk(reg_896__clk),
    .in(reg_896__in),
    .out(reg_896__out)
  );

  //Wire declarations for instance 'reg_897' (Module coreir_reg)
  wire  reg_897__clk;
  wire [15:0] reg_897__in;
  wire [15:0] reg_897__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_897(
    .clk(reg_897__clk),
    .in(reg_897__in),
    .out(reg_897__out)
  );

  //Wire declarations for instance 'reg_898' (Module coreir_reg)
  wire  reg_898__clk;
  wire [15:0] reg_898__in;
  wire [15:0] reg_898__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_898(
    .clk(reg_898__clk),
    .in(reg_898__in),
    .out(reg_898__out)
  );

  //Wire declarations for instance 'reg_899' (Module coreir_reg)
  wire  reg_899__clk;
  wire [15:0] reg_899__in;
  wire [15:0] reg_899__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_899(
    .clk(reg_899__clk),
    .in(reg_899__in),
    .out(reg_899__out)
  );

  //Wire declarations for instance 'reg_9' (Module coreir_reg)
  wire  reg_9__clk;
  wire [15:0] reg_9__in;
  wire [15:0] reg_9__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_9(
    .clk(reg_9__clk),
    .in(reg_9__in),
    .out(reg_9__out)
  );

  //Wire declarations for instance 'reg_90' (Module coreir_reg)
  wire  reg_90__clk;
  wire [15:0] reg_90__in;
  wire [15:0] reg_90__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_90(
    .clk(reg_90__clk),
    .in(reg_90__in),
    .out(reg_90__out)
  );

  //Wire declarations for instance 'reg_900' (Module coreir_reg)
  wire  reg_900__clk;
  wire [15:0] reg_900__in;
  wire [15:0] reg_900__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_900(
    .clk(reg_900__clk),
    .in(reg_900__in),
    .out(reg_900__out)
  );

  //Wire declarations for instance 'reg_901' (Module coreir_reg)
  wire  reg_901__clk;
  wire [15:0] reg_901__in;
  wire [15:0] reg_901__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_901(
    .clk(reg_901__clk),
    .in(reg_901__in),
    .out(reg_901__out)
  );

  //Wire declarations for instance 'reg_902' (Module coreir_reg)
  wire  reg_902__clk;
  wire [15:0] reg_902__in;
  wire [15:0] reg_902__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_902(
    .clk(reg_902__clk),
    .in(reg_902__in),
    .out(reg_902__out)
  );

  //Wire declarations for instance 'reg_903' (Module coreir_reg)
  wire  reg_903__clk;
  wire [15:0] reg_903__in;
  wire [15:0] reg_903__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_903(
    .clk(reg_903__clk),
    .in(reg_903__in),
    .out(reg_903__out)
  );

  //Wire declarations for instance 'reg_904' (Module coreir_reg)
  wire  reg_904__clk;
  wire [15:0] reg_904__in;
  wire [15:0] reg_904__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_904(
    .clk(reg_904__clk),
    .in(reg_904__in),
    .out(reg_904__out)
  );

  //Wire declarations for instance 'reg_905' (Module coreir_reg)
  wire  reg_905__clk;
  wire [15:0] reg_905__in;
  wire [15:0] reg_905__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_905(
    .clk(reg_905__clk),
    .in(reg_905__in),
    .out(reg_905__out)
  );

  //Wire declarations for instance 'reg_906' (Module coreir_reg)
  wire  reg_906__clk;
  wire [15:0] reg_906__in;
  wire [15:0] reg_906__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_906(
    .clk(reg_906__clk),
    .in(reg_906__in),
    .out(reg_906__out)
  );

  //Wire declarations for instance 'reg_907' (Module coreir_reg)
  wire  reg_907__clk;
  wire [15:0] reg_907__in;
  wire [15:0] reg_907__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_907(
    .clk(reg_907__clk),
    .in(reg_907__in),
    .out(reg_907__out)
  );

  //Wire declarations for instance 'reg_908' (Module coreir_reg)
  wire  reg_908__clk;
  wire [15:0] reg_908__in;
  wire [15:0] reg_908__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_908(
    .clk(reg_908__clk),
    .in(reg_908__in),
    .out(reg_908__out)
  );

  //Wire declarations for instance 'reg_909' (Module coreir_reg)
  wire  reg_909__clk;
  wire [15:0] reg_909__in;
  wire [15:0] reg_909__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_909(
    .clk(reg_909__clk),
    .in(reg_909__in),
    .out(reg_909__out)
  );

  //Wire declarations for instance 'reg_91' (Module coreir_reg)
  wire  reg_91__clk;
  wire [15:0] reg_91__in;
  wire [15:0] reg_91__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_91(
    .clk(reg_91__clk),
    .in(reg_91__in),
    .out(reg_91__out)
  );

  //Wire declarations for instance 'reg_910' (Module coreir_reg)
  wire  reg_910__clk;
  wire [15:0] reg_910__in;
  wire [15:0] reg_910__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_910(
    .clk(reg_910__clk),
    .in(reg_910__in),
    .out(reg_910__out)
  );

  //Wire declarations for instance 'reg_911' (Module coreir_reg)
  wire  reg_911__clk;
  wire [15:0] reg_911__in;
  wire [15:0] reg_911__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_911(
    .clk(reg_911__clk),
    .in(reg_911__in),
    .out(reg_911__out)
  );

  //Wire declarations for instance 'reg_912' (Module coreir_reg)
  wire  reg_912__clk;
  wire [15:0] reg_912__in;
  wire [15:0] reg_912__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_912(
    .clk(reg_912__clk),
    .in(reg_912__in),
    .out(reg_912__out)
  );

  //Wire declarations for instance 'reg_913' (Module coreir_reg)
  wire  reg_913__clk;
  wire [15:0] reg_913__in;
  wire [15:0] reg_913__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_913(
    .clk(reg_913__clk),
    .in(reg_913__in),
    .out(reg_913__out)
  );

  //Wire declarations for instance 'reg_914' (Module coreir_reg)
  wire  reg_914__clk;
  wire [15:0] reg_914__in;
  wire [15:0] reg_914__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_914(
    .clk(reg_914__clk),
    .in(reg_914__in),
    .out(reg_914__out)
  );

  //Wire declarations for instance 'reg_915' (Module coreir_reg)
  wire  reg_915__clk;
  wire [15:0] reg_915__in;
  wire [15:0] reg_915__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_915(
    .clk(reg_915__clk),
    .in(reg_915__in),
    .out(reg_915__out)
  );

  //Wire declarations for instance 'reg_916' (Module coreir_reg)
  wire  reg_916__clk;
  wire [15:0] reg_916__in;
  wire [15:0] reg_916__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_916(
    .clk(reg_916__clk),
    .in(reg_916__in),
    .out(reg_916__out)
  );

  //Wire declarations for instance 'reg_917' (Module coreir_reg)
  wire  reg_917__clk;
  wire [15:0] reg_917__in;
  wire [15:0] reg_917__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_917(
    .clk(reg_917__clk),
    .in(reg_917__in),
    .out(reg_917__out)
  );

  //Wire declarations for instance 'reg_918' (Module coreir_reg)
  wire  reg_918__clk;
  wire [15:0] reg_918__in;
  wire [15:0] reg_918__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_918(
    .clk(reg_918__clk),
    .in(reg_918__in),
    .out(reg_918__out)
  );

  //Wire declarations for instance 'reg_919' (Module coreir_reg)
  wire  reg_919__clk;
  wire [15:0] reg_919__in;
  wire [15:0] reg_919__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_919(
    .clk(reg_919__clk),
    .in(reg_919__in),
    .out(reg_919__out)
  );

  //Wire declarations for instance 'reg_92' (Module coreir_reg)
  wire  reg_92__clk;
  wire [15:0] reg_92__in;
  wire [15:0] reg_92__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_92(
    .clk(reg_92__clk),
    .in(reg_92__in),
    .out(reg_92__out)
  );

  //Wire declarations for instance 'reg_920' (Module coreir_reg)
  wire  reg_920__clk;
  wire [15:0] reg_920__in;
  wire [15:0] reg_920__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_920(
    .clk(reg_920__clk),
    .in(reg_920__in),
    .out(reg_920__out)
  );

  //Wire declarations for instance 'reg_921' (Module coreir_reg)
  wire  reg_921__clk;
  wire [15:0] reg_921__in;
  wire [15:0] reg_921__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_921(
    .clk(reg_921__clk),
    .in(reg_921__in),
    .out(reg_921__out)
  );

  //Wire declarations for instance 'reg_922' (Module coreir_reg)
  wire  reg_922__clk;
  wire [15:0] reg_922__in;
  wire [15:0] reg_922__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_922(
    .clk(reg_922__clk),
    .in(reg_922__in),
    .out(reg_922__out)
  );

  //Wire declarations for instance 'reg_923' (Module coreir_reg)
  wire  reg_923__clk;
  wire [15:0] reg_923__in;
  wire [15:0] reg_923__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_923(
    .clk(reg_923__clk),
    .in(reg_923__in),
    .out(reg_923__out)
  );

  //Wire declarations for instance 'reg_924' (Module coreir_reg)
  wire  reg_924__clk;
  wire [15:0] reg_924__in;
  wire [15:0] reg_924__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_924(
    .clk(reg_924__clk),
    .in(reg_924__in),
    .out(reg_924__out)
  );

  //Wire declarations for instance 'reg_925' (Module coreir_reg)
  wire  reg_925__clk;
  wire [15:0] reg_925__in;
  wire [15:0] reg_925__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_925(
    .clk(reg_925__clk),
    .in(reg_925__in),
    .out(reg_925__out)
  );

  //Wire declarations for instance 'reg_926' (Module coreir_reg)
  wire  reg_926__clk;
  wire [15:0] reg_926__in;
  wire [15:0] reg_926__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_926(
    .clk(reg_926__clk),
    .in(reg_926__in),
    .out(reg_926__out)
  );

  //Wire declarations for instance 'reg_927' (Module coreir_reg)
  wire  reg_927__clk;
  wire [15:0] reg_927__in;
  wire [15:0] reg_927__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_927(
    .clk(reg_927__clk),
    .in(reg_927__in),
    .out(reg_927__out)
  );

  //Wire declarations for instance 'reg_928' (Module coreir_reg)
  wire  reg_928__clk;
  wire [15:0] reg_928__in;
  wire [15:0] reg_928__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_928(
    .clk(reg_928__clk),
    .in(reg_928__in),
    .out(reg_928__out)
  );

  //Wire declarations for instance 'reg_929' (Module coreir_reg)
  wire  reg_929__clk;
  wire [15:0] reg_929__in;
  wire [15:0] reg_929__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_929(
    .clk(reg_929__clk),
    .in(reg_929__in),
    .out(reg_929__out)
  );

  //Wire declarations for instance 'reg_93' (Module coreir_reg)
  wire  reg_93__clk;
  wire [15:0] reg_93__in;
  wire [15:0] reg_93__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_93(
    .clk(reg_93__clk),
    .in(reg_93__in),
    .out(reg_93__out)
  );

  //Wire declarations for instance 'reg_930' (Module coreir_reg)
  wire  reg_930__clk;
  wire [15:0] reg_930__in;
  wire [15:0] reg_930__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_930(
    .clk(reg_930__clk),
    .in(reg_930__in),
    .out(reg_930__out)
  );

  //Wire declarations for instance 'reg_931' (Module coreir_reg)
  wire  reg_931__clk;
  wire [15:0] reg_931__in;
  wire [15:0] reg_931__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_931(
    .clk(reg_931__clk),
    .in(reg_931__in),
    .out(reg_931__out)
  );

  //Wire declarations for instance 'reg_932' (Module coreir_reg)
  wire  reg_932__clk;
  wire [15:0] reg_932__in;
  wire [15:0] reg_932__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_932(
    .clk(reg_932__clk),
    .in(reg_932__in),
    .out(reg_932__out)
  );

  //Wire declarations for instance 'reg_933' (Module coreir_reg)
  wire  reg_933__clk;
  wire [15:0] reg_933__in;
  wire [15:0] reg_933__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_933(
    .clk(reg_933__clk),
    .in(reg_933__in),
    .out(reg_933__out)
  );

  //Wire declarations for instance 'reg_934' (Module coreir_reg)
  wire  reg_934__clk;
  wire [15:0] reg_934__in;
  wire [15:0] reg_934__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_934(
    .clk(reg_934__clk),
    .in(reg_934__in),
    .out(reg_934__out)
  );

  //Wire declarations for instance 'reg_935' (Module coreir_reg)
  wire  reg_935__clk;
  wire [15:0] reg_935__in;
  wire [15:0] reg_935__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_935(
    .clk(reg_935__clk),
    .in(reg_935__in),
    .out(reg_935__out)
  );

  //Wire declarations for instance 'reg_936' (Module coreir_reg)
  wire  reg_936__clk;
  wire [15:0] reg_936__in;
  wire [15:0] reg_936__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_936(
    .clk(reg_936__clk),
    .in(reg_936__in),
    .out(reg_936__out)
  );

  //Wire declarations for instance 'reg_937' (Module coreir_reg)
  wire  reg_937__clk;
  wire [15:0] reg_937__in;
  wire [15:0] reg_937__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_937(
    .clk(reg_937__clk),
    .in(reg_937__in),
    .out(reg_937__out)
  );

  //Wire declarations for instance 'reg_938' (Module coreir_reg)
  wire  reg_938__clk;
  wire [15:0] reg_938__in;
  wire [15:0] reg_938__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_938(
    .clk(reg_938__clk),
    .in(reg_938__in),
    .out(reg_938__out)
  );

  //Wire declarations for instance 'reg_939' (Module coreir_reg)
  wire  reg_939__clk;
  wire [15:0] reg_939__in;
  wire [15:0] reg_939__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_939(
    .clk(reg_939__clk),
    .in(reg_939__in),
    .out(reg_939__out)
  );

  //Wire declarations for instance 'reg_94' (Module coreir_reg)
  wire  reg_94__clk;
  wire [15:0] reg_94__in;
  wire [15:0] reg_94__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_94(
    .clk(reg_94__clk),
    .in(reg_94__in),
    .out(reg_94__out)
  );

  //Wire declarations for instance 'reg_940' (Module coreir_reg)
  wire  reg_940__clk;
  wire [15:0] reg_940__in;
  wire [15:0] reg_940__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_940(
    .clk(reg_940__clk),
    .in(reg_940__in),
    .out(reg_940__out)
  );

  //Wire declarations for instance 'reg_941' (Module coreir_reg)
  wire  reg_941__clk;
  wire [15:0] reg_941__in;
  wire [15:0] reg_941__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_941(
    .clk(reg_941__clk),
    .in(reg_941__in),
    .out(reg_941__out)
  );

  //Wire declarations for instance 'reg_942' (Module coreir_reg)
  wire  reg_942__clk;
  wire [15:0] reg_942__in;
  wire [15:0] reg_942__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_942(
    .clk(reg_942__clk),
    .in(reg_942__in),
    .out(reg_942__out)
  );

  //Wire declarations for instance 'reg_943' (Module coreir_reg)
  wire  reg_943__clk;
  wire [15:0] reg_943__in;
  wire [15:0] reg_943__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_943(
    .clk(reg_943__clk),
    .in(reg_943__in),
    .out(reg_943__out)
  );

  //Wire declarations for instance 'reg_944' (Module coreir_reg)
  wire  reg_944__clk;
  wire [15:0] reg_944__in;
  wire [15:0] reg_944__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_944(
    .clk(reg_944__clk),
    .in(reg_944__in),
    .out(reg_944__out)
  );

  //Wire declarations for instance 'reg_945' (Module coreir_reg)
  wire  reg_945__clk;
  wire [15:0] reg_945__in;
  wire [15:0] reg_945__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_945(
    .clk(reg_945__clk),
    .in(reg_945__in),
    .out(reg_945__out)
  );

  //Wire declarations for instance 'reg_946' (Module coreir_reg)
  wire  reg_946__clk;
  wire [15:0] reg_946__in;
  wire [15:0] reg_946__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_946(
    .clk(reg_946__clk),
    .in(reg_946__in),
    .out(reg_946__out)
  );

  //Wire declarations for instance 'reg_947' (Module coreir_reg)
  wire  reg_947__clk;
  wire [15:0] reg_947__in;
  wire [15:0] reg_947__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_947(
    .clk(reg_947__clk),
    .in(reg_947__in),
    .out(reg_947__out)
  );

  //Wire declarations for instance 'reg_948' (Module coreir_reg)
  wire  reg_948__clk;
  wire [15:0] reg_948__in;
  wire [15:0] reg_948__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_948(
    .clk(reg_948__clk),
    .in(reg_948__in),
    .out(reg_948__out)
  );

  //Wire declarations for instance 'reg_949' (Module coreir_reg)
  wire  reg_949__clk;
  wire [15:0] reg_949__in;
  wire [15:0] reg_949__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_949(
    .clk(reg_949__clk),
    .in(reg_949__in),
    .out(reg_949__out)
  );

  //Wire declarations for instance 'reg_95' (Module coreir_reg)
  wire  reg_95__clk;
  wire [15:0] reg_95__in;
  wire [15:0] reg_95__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_95(
    .clk(reg_95__clk),
    .in(reg_95__in),
    .out(reg_95__out)
  );

  //Wire declarations for instance 'reg_950' (Module coreir_reg)
  wire  reg_950__clk;
  wire [15:0] reg_950__in;
  wire [15:0] reg_950__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_950(
    .clk(reg_950__clk),
    .in(reg_950__in),
    .out(reg_950__out)
  );

  //Wire declarations for instance 'reg_951' (Module coreir_reg)
  wire  reg_951__clk;
  wire [15:0] reg_951__in;
  wire [15:0] reg_951__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_951(
    .clk(reg_951__clk),
    .in(reg_951__in),
    .out(reg_951__out)
  );

  //Wire declarations for instance 'reg_952' (Module coreir_reg)
  wire  reg_952__clk;
  wire [15:0] reg_952__in;
  wire [15:0] reg_952__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_952(
    .clk(reg_952__clk),
    .in(reg_952__in),
    .out(reg_952__out)
  );

  //Wire declarations for instance 'reg_953' (Module coreir_reg)
  wire  reg_953__clk;
  wire [15:0] reg_953__in;
  wire [15:0] reg_953__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_953(
    .clk(reg_953__clk),
    .in(reg_953__in),
    .out(reg_953__out)
  );

  //Wire declarations for instance 'reg_954' (Module coreir_reg)
  wire  reg_954__clk;
  wire [15:0] reg_954__in;
  wire [15:0] reg_954__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_954(
    .clk(reg_954__clk),
    .in(reg_954__in),
    .out(reg_954__out)
  );

  //Wire declarations for instance 'reg_955' (Module coreir_reg)
  wire  reg_955__clk;
  wire [15:0] reg_955__in;
  wire [15:0] reg_955__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_955(
    .clk(reg_955__clk),
    .in(reg_955__in),
    .out(reg_955__out)
  );

  //Wire declarations for instance 'reg_956' (Module coreir_reg)
  wire  reg_956__clk;
  wire [15:0] reg_956__in;
  wire [15:0] reg_956__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_956(
    .clk(reg_956__clk),
    .in(reg_956__in),
    .out(reg_956__out)
  );

  //Wire declarations for instance 'reg_957' (Module coreir_reg)
  wire  reg_957__clk;
  wire [15:0] reg_957__in;
  wire [15:0] reg_957__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_957(
    .clk(reg_957__clk),
    .in(reg_957__in),
    .out(reg_957__out)
  );

  //Wire declarations for instance 'reg_958' (Module coreir_reg)
  wire  reg_958__clk;
  wire [15:0] reg_958__in;
  wire [15:0] reg_958__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_958(
    .clk(reg_958__clk),
    .in(reg_958__in),
    .out(reg_958__out)
  );

  //Wire declarations for instance 'reg_959' (Module coreir_reg)
  wire  reg_959__clk;
  wire [15:0] reg_959__in;
  wire [15:0] reg_959__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_959(
    .clk(reg_959__clk),
    .in(reg_959__in),
    .out(reg_959__out)
  );

  //Wire declarations for instance 'reg_96' (Module coreir_reg)
  wire  reg_96__clk;
  wire [15:0] reg_96__in;
  wire [15:0] reg_96__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_96(
    .clk(reg_96__clk),
    .in(reg_96__in),
    .out(reg_96__out)
  );

  //Wire declarations for instance 'reg_960' (Module coreir_reg)
  wire  reg_960__clk;
  wire [15:0] reg_960__in;
  wire [15:0] reg_960__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_960(
    .clk(reg_960__clk),
    .in(reg_960__in),
    .out(reg_960__out)
  );

  //Wire declarations for instance 'reg_961' (Module coreir_reg)
  wire  reg_961__clk;
  wire [15:0] reg_961__in;
  wire [15:0] reg_961__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_961(
    .clk(reg_961__clk),
    .in(reg_961__in),
    .out(reg_961__out)
  );

  //Wire declarations for instance 'reg_962' (Module coreir_reg)
  wire  reg_962__clk;
  wire [15:0] reg_962__in;
  wire [15:0] reg_962__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_962(
    .clk(reg_962__clk),
    .in(reg_962__in),
    .out(reg_962__out)
  );

  //Wire declarations for instance 'reg_963' (Module coreir_reg)
  wire  reg_963__clk;
  wire [15:0] reg_963__in;
  wire [15:0] reg_963__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_963(
    .clk(reg_963__clk),
    .in(reg_963__in),
    .out(reg_963__out)
  );

  //Wire declarations for instance 'reg_964' (Module coreir_reg)
  wire  reg_964__clk;
  wire [15:0] reg_964__in;
  wire [15:0] reg_964__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_964(
    .clk(reg_964__clk),
    .in(reg_964__in),
    .out(reg_964__out)
  );

  //Wire declarations for instance 'reg_965' (Module coreir_reg)
  wire  reg_965__clk;
  wire [15:0] reg_965__in;
  wire [15:0] reg_965__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_965(
    .clk(reg_965__clk),
    .in(reg_965__in),
    .out(reg_965__out)
  );

  //Wire declarations for instance 'reg_966' (Module coreir_reg)
  wire  reg_966__clk;
  wire [15:0] reg_966__in;
  wire [15:0] reg_966__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_966(
    .clk(reg_966__clk),
    .in(reg_966__in),
    .out(reg_966__out)
  );

  //Wire declarations for instance 'reg_967' (Module coreir_reg)
  wire  reg_967__clk;
  wire [15:0] reg_967__in;
  wire [15:0] reg_967__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_967(
    .clk(reg_967__clk),
    .in(reg_967__in),
    .out(reg_967__out)
  );

  //Wire declarations for instance 'reg_968' (Module coreir_reg)
  wire  reg_968__clk;
  wire [15:0] reg_968__in;
  wire [15:0] reg_968__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_968(
    .clk(reg_968__clk),
    .in(reg_968__in),
    .out(reg_968__out)
  );

  //Wire declarations for instance 'reg_969' (Module coreir_reg)
  wire  reg_969__clk;
  wire [15:0] reg_969__in;
  wire [15:0] reg_969__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_969(
    .clk(reg_969__clk),
    .in(reg_969__in),
    .out(reg_969__out)
  );

  //Wire declarations for instance 'reg_97' (Module coreir_reg)
  wire  reg_97__clk;
  wire [15:0] reg_97__in;
  wire [15:0] reg_97__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_97(
    .clk(reg_97__clk),
    .in(reg_97__in),
    .out(reg_97__out)
  );

  //Wire declarations for instance 'reg_970' (Module coreir_reg)
  wire  reg_970__clk;
  wire [15:0] reg_970__in;
  wire [15:0] reg_970__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_970(
    .clk(reg_970__clk),
    .in(reg_970__in),
    .out(reg_970__out)
  );

  //Wire declarations for instance 'reg_971' (Module coreir_reg)
  wire  reg_971__clk;
  wire [15:0] reg_971__in;
  wire [15:0] reg_971__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_971(
    .clk(reg_971__clk),
    .in(reg_971__in),
    .out(reg_971__out)
  );

  //Wire declarations for instance 'reg_972' (Module coreir_reg)
  wire  reg_972__clk;
  wire [15:0] reg_972__in;
  wire [15:0] reg_972__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_972(
    .clk(reg_972__clk),
    .in(reg_972__in),
    .out(reg_972__out)
  );

  //Wire declarations for instance 'reg_973' (Module coreir_reg)
  wire  reg_973__clk;
  wire [15:0] reg_973__in;
  wire [15:0] reg_973__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_973(
    .clk(reg_973__clk),
    .in(reg_973__in),
    .out(reg_973__out)
  );

  //Wire declarations for instance 'reg_974' (Module coreir_reg)
  wire  reg_974__clk;
  wire [15:0] reg_974__in;
  wire [15:0] reg_974__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_974(
    .clk(reg_974__clk),
    .in(reg_974__in),
    .out(reg_974__out)
  );

  //Wire declarations for instance 'reg_975' (Module coreir_reg)
  wire  reg_975__clk;
  wire [15:0] reg_975__in;
  wire [15:0] reg_975__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_975(
    .clk(reg_975__clk),
    .in(reg_975__in),
    .out(reg_975__out)
  );

  //Wire declarations for instance 'reg_976' (Module coreir_reg)
  wire  reg_976__clk;
  wire [15:0] reg_976__in;
  wire [15:0] reg_976__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_976(
    .clk(reg_976__clk),
    .in(reg_976__in),
    .out(reg_976__out)
  );

  //Wire declarations for instance 'reg_977' (Module coreir_reg)
  wire  reg_977__clk;
  wire [15:0] reg_977__in;
  wire [15:0] reg_977__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_977(
    .clk(reg_977__clk),
    .in(reg_977__in),
    .out(reg_977__out)
  );

  //Wire declarations for instance 'reg_978' (Module coreir_reg)
  wire  reg_978__clk;
  wire [15:0] reg_978__in;
  wire [15:0] reg_978__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_978(
    .clk(reg_978__clk),
    .in(reg_978__in),
    .out(reg_978__out)
  );

  //Wire declarations for instance 'reg_979' (Module coreir_reg)
  wire  reg_979__clk;
  wire [15:0] reg_979__in;
  wire [15:0] reg_979__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_979(
    .clk(reg_979__clk),
    .in(reg_979__in),
    .out(reg_979__out)
  );

  //Wire declarations for instance 'reg_98' (Module coreir_reg)
  wire  reg_98__clk;
  wire [15:0] reg_98__in;
  wire [15:0] reg_98__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_98(
    .clk(reg_98__clk),
    .in(reg_98__in),
    .out(reg_98__out)
  );

  //Wire declarations for instance 'reg_980' (Module coreir_reg)
  wire  reg_980__clk;
  wire [15:0] reg_980__in;
  wire [15:0] reg_980__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_980(
    .clk(reg_980__clk),
    .in(reg_980__in),
    .out(reg_980__out)
  );

  //Wire declarations for instance 'reg_981' (Module coreir_reg)
  wire  reg_981__clk;
  wire [15:0] reg_981__in;
  wire [15:0] reg_981__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_981(
    .clk(reg_981__clk),
    .in(reg_981__in),
    .out(reg_981__out)
  );

  //Wire declarations for instance 'reg_982' (Module coreir_reg)
  wire  reg_982__clk;
  wire [15:0] reg_982__in;
  wire [15:0] reg_982__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_982(
    .clk(reg_982__clk),
    .in(reg_982__in),
    .out(reg_982__out)
  );

  //Wire declarations for instance 'reg_983' (Module coreir_reg)
  wire  reg_983__clk;
  wire [15:0] reg_983__in;
  wire [15:0] reg_983__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_983(
    .clk(reg_983__clk),
    .in(reg_983__in),
    .out(reg_983__out)
  );

  //Wire declarations for instance 'reg_984' (Module coreir_reg)
  wire  reg_984__clk;
  wire [15:0] reg_984__in;
  wire [15:0] reg_984__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_984(
    .clk(reg_984__clk),
    .in(reg_984__in),
    .out(reg_984__out)
  );

  //Wire declarations for instance 'reg_985' (Module coreir_reg)
  wire  reg_985__clk;
  wire [15:0] reg_985__in;
  wire [15:0] reg_985__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_985(
    .clk(reg_985__clk),
    .in(reg_985__in),
    .out(reg_985__out)
  );

  //Wire declarations for instance 'reg_986' (Module coreir_reg)
  wire  reg_986__clk;
  wire [15:0] reg_986__in;
  wire [15:0] reg_986__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_986(
    .clk(reg_986__clk),
    .in(reg_986__in),
    .out(reg_986__out)
  );

  //Wire declarations for instance 'reg_987' (Module coreir_reg)
  wire  reg_987__clk;
  wire [15:0] reg_987__in;
  wire [15:0] reg_987__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_987(
    .clk(reg_987__clk),
    .in(reg_987__in),
    .out(reg_987__out)
  );

  //Wire declarations for instance 'reg_988' (Module coreir_reg)
  wire  reg_988__clk;
  wire [15:0] reg_988__in;
  wire [15:0] reg_988__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_988(
    .clk(reg_988__clk),
    .in(reg_988__in),
    .out(reg_988__out)
  );

  //Wire declarations for instance 'reg_989' (Module coreir_reg)
  wire  reg_989__clk;
  wire [15:0] reg_989__in;
  wire [15:0] reg_989__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_989(
    .clk(reg_989__clk),
    .in(reg_989__in),
    .out(reg_989__out)
  );

  //Wire declarations for instance 'reg_99' (Module coreir_reg)
  wire  reg_99__clk;
  wire [15:0] reg_99__in;
  wire [15:0] reg_99__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_99(
    .clk(reg_99__clk),
    .in(reg_99__in),
    .out(reg_99__out)
  );

  //Wire declarations for instance 'reg_990' (Module coreir_reg)
  wire  reg_990__clk;
  wire [15:0] reg_990__in;
  wire [15:0] reg_990__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_990(
    .clk(reg_990__clk),
    .in(reg_990__in),
    .out(reg_990__out)
  );

  //Wire declarations for instance 'reg_991' (Module coreir_reg)
  wire  reg_991__clk;
  wire [15:0] reg_991__in;
  wire [15:0] reg_991__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_991(
    .clk(reg_991__clk),
    .in(reg_991__in),
    .out(reg_991__out)
  );

  //Wire declarations for instance 'reg_992' (Module coreir_reg)
  wire  reg_992__clk;
  wire [15:0] reg_992__in;
  wire [15:0] reg_992__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_992(
    .clk(reg_992__clk),
    .in(reg_992__in),
    .out(reg_992__out)
  );

  //Wire declarations for instance 'reg_993' (Module coreir_reg)
  wire  reg_993__clk;
  wire [15:0] reg_993__in;
  wire [15:0] reg_993__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_993(
    .clk(reg_993__clk),
    .in(reg_993__in),
    .out(reg_993__out)
  );

  //Wire declarations for instance 'reg_994' (Module coreir_reg)
  wire  reg_994__clk;
  wire [15:0] reg_994__in;
  wire [15:0] reg_994__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_994(
    .clk(reg_994__clk),
    .in(reg_994__in),
    .out(reg_994__out)
  );

  //Wire declarations for instance 'reg_995' (Module coreir_reg)
  wire  reg_995__clk;
  wire [15:0] reg_995__in;
  wire [15:0] reg_995__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_995(
    .clk(reg_995__clk),
    .in(reg_995__in),
    .out(reg_995__out)
  );

  //Wire declarations for instance 'reg_996' (Module coreir_reg)
  wire  reg_996__clk;
  wire [15:0] reg_996__in;
  wire [15:0] reg_996__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_996(
    .clk(reg_996__clk),
    .in(reg_996__in),
    .out(reg_996__out)
  );

  //Wire declarations for instance 'reg_997' (Module coreir_reg)
  wire  reg_997__clk;
  wire [15:0] reg_997__in;
  wire [15:0] reg_997__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_997(
    .clk(reg_997__clk),
    .in(reg_997__in),
    .out(reg_997__out)
  );

  //Wire declarations for instance 'reg_998' (Module coreir_reg)
  wire  reg_998__clk;
  wire [15:0] reg_998__in;
  wire [15:0] reg_998__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_998(
    .clk(reg_998__clk),
    .in(reg_998__in),
    .out(reg_998__out)
  );

  //Wire declarations for instance 'reg_999' (Module coreir_reg)
  wire  reg_999__clk;
  wire [15:0] reg_999__in;
  wire [15:0] reg_999__out;
  coreir_reg #(.init(16'd0),.width(16)) reg_999(
    .clk(reg_999__clk),
    .in(reg_999__in),
    .out(reg_999__out)
  );

  //All the connections
  assign and_0__in0[15:0] = in_0[15:0];
  assign and_0__in1[15:0] = in_1[15:0];
  assign reg_0__in[15:0] = and_0__out[15:0];
  assign and_10__in0[15:0] = in_20[15:0];
  assign and_10__in1[15:0] = in_21[15:0];
  assign reg_10__in[15:0] = and_10__out[15:0];
  assign and_100__in0[15:0] = in_200[15:0];
  assign and_100__in1[15:0] = in_201[15:0];
  assign reg_100__in[15:0] = and_100__out[15:0];
  assign and_102__in0[15:0] = in_204[15:0];
  assign and_102__in1[15:0] = in_205[15:0];
  assign reg_102__in[15:0] = and_102__out[15:0];
  assign and_104__in0[15:0] = in_208[15:0];
  assign and_104__in1[15:0] = in_209[15:0];
  assign reg_104__in[15:0] = and_104__out[15:0];
  assign and_106__in0[15:0] = in_212[15:0];
  assign and_106__in1[15:0] = in_213[15:0];
  assign reg_106__in[15:0] = and_106__out[15:0];
  assign and_108__in0[15:0] = in_216[15:0];
  assign and_108__in1[15:0] = in_217[15:0];
  assign reg_108__in[15:0] = and_108__out[15:0];
  assign and_110__in0[15:0] = in_220[15:0];
  assign and_110__in1[15:0] = in_221[15:0];
  assign reg_110__in[15:0] = and_110__out[15:0];
  assign and_112__in0[15:0] = in_224[15:0];
  assign and_112__in1[15:0] = in_225[15:0];
  assign reg_112__in[15:0] = and_112__out[15:0];
  assign and_114__in0[15:0] = in_228[15:0];
  assign and_114__in1[15:0] = in_229[15:0];
  assign reg_114__in[15:0] = and_114__out[15:0];
  assign and_116__in0[15:0] = in_232[15:0];
  assign and_116__in1[15:0] = in_233[15:0];
  assign reg_116__in[15:0] = and_116__out[15:0];
  assign and_118__in0[15:0] = in_236[15:0];
  assign and_118__in1[15:0] = in_237[15:0];
  assign reg_118__in[15:0] = and_118__out[15:0];
  assign and_12__in0[15:0] = in_24[15:0];
  assign and_12__in1[15:0] = in_25[15:0];
  assign reg_12__in[15:0] = and_12__out[15:0];
  assign and_120__in0[15:0] = in_240[15:0];
  assign and_120__in1[15:0] = in_241[15:0];
  assign reg_120__in[15:0] = and_120__out[15:0];
  assign and_122__in0[15:0] = in_244[15:0];
  assign and_122__in1[15:0] = in_245[15:0];
  assign reg_122__in[15:0] = and_122__out[15:0];
  assign and_124__in0[15:0] = in_248[15:0];
  assign and_124__in1[15:0] = in_249[15:0];
  assign reg_124__in[15:0] = and_124__out[15:0];
  assign and_126__in0[15:0] = in_252[15:0];
  assign and_126__in1[15:0] = in_253[15:0];
  assign reg_126__in[15:0] = and_126__out[15:0];
  assign and_128__in0[15:0] = in_256[15:0];
  assign and_128__in1[15:0] = in_257[15:0];
  assign reg_128__in[15:0] = and_128__out[15:0];
  assign and_130__in0[15:0] = in_260[15:0];
  assign and_130__in1[15:0] = in_261[15:0];
  assign reg_130__in[15:0] = and_130__out[15:0];
  assign and_132__in0[15:0] = in_264[15:0];
  assign and_132__in1[15:0] = in_265[15:0];
  assign reg_132__in[15:0] = and_132__out[15:0];
  assign and_134__in0[15:0] = in_268[15:0];
  assign and_134__in1[15:0] = in_269[15:0];
  assign reg_134__in[15:0] = and_134__out[15:0];
  assign and_136__in0[15:0] = in_272[15:0];
  assign and_136__in1[15:0] = in_273[15:0];
  assign reg_136__in[15:0] = and_136__out[15:0];
  assign and_138__in0[15:0] = in_276[15:0];
  assign and_138__in1[15:0] = in_277[15:0];
  assign reg_138__in[15:0] = and_138__out[15:0];
  assign and_14__in0[15:0] = in_28[15:0];
  assign and_14__in1[15:0] = in_29[15:0];
  assign reg_14__in[15:0] = and_14__out[15:0];
  assign and_140__in0[15:0] = in_280[15:0];
  assign and_140__in1[15:0] = in_281[15:0];
  assign reg_140__in[15:0] = and_140__out[15:0];
  assign and_142__in0[15:0] = in_284[15:0];
  assign and_142__in1[15:0] = in_285[15:0];
  assign reg_142__in[15:0] = and_142__out[15:0];
  assign and_144__in0[15:0] = in_288[15:0];
  assign and_144__in1[15:0] = in_289[15:0];
  assign reg_144__in[15:0] = and_144__out[15:0];
  assign and_146__in0[15:0] = in_292[15:0];
  assign and_146__in1[15:0] = in_293[15:0];
  assign reg_146__in[15:0] = and_146__out[15:0];
  assign and_148__in0[15:0] = in_296[15:0];
  assign and_148__in1[15:0] = in_297[15:0];
  assign reg_148__in[15:0] = and_148__out[15:0];
  assign and_150__in0[15:0] = in_300[15:0];
  assign and_150__in1[15:0] = in_301[15:0];
  assign reg_150__in[15:0] = and_150__out[15:0];
  assign and_152__in0[15:0] = in_304[15:0];
  assign and_152__in1[15:0] = in_305[15:0];
  assign reg_152__in[15:0] = and_152__out[15:0];
  assign and_154__in0[15:0] = in_308[15:0];
  assign and_154__in1[15:0] = in_309[15:0];
  assign reg_154__in[15:0] = and_154__out[15:0];
  assign and_156__in0[15:0] = in_312[15:0];
  assign and_156__in1[15:0] = in_313[15:0];
  assign reg_156__in[15:0] = and_156__out[15:0];
  assign and_158__in0[15:0] = in_316[15:0];
  assign and_158__in1[15:0] = in_317[15:0];
  assign reg_158__in[15:0] = and_158__out[15:0];
  assign and_16__in0[15:0] = in_32[15:0];
  assign and_16__in1[15:0] = in_33[15:0];
  assign reg_16__in[15:0] = and_16__out[15:0];
  assign and_160__in0[15:0] = in_320[15:0];
  assign and_160__in1[15:0] = in_321[15:0];
  assign reg_160__in[15:0] = and_160__out[15:0];
  assign and_162__in0[15:0] = in_324[15:0];
  assign and_162__in1[15:0] = in_325[15:0];
  assign reg_162__in[15:0] = and_162__out[15:0];
  assign and_164__in0[15:0] = in_328[15:0];
  assign and_164__in1[15:0] = in_329[15:0];
  assign reg_164__in[15:0] = and_164__out[15:0];
  assign and_166__in0[15:0] = in_332[15:0];
  assign and_166__in1[15:0] = in_333[15:0];
  assign reg_166__in[15:0] = and_166__out[15:0];
  assign and_168__in0[15:0] = in_336[15:0];
  assign and_168__in1[15:0] = in_337[15:0];
  assign reg_168__in[15:0] = and_168__out[15:0];
  assign and_170__in0[15:0] = in_340[15:0];
  assign and_170__in1[15:0] = in_341[15:0];
  assign reg_170__in[15:0] = and_170__out[15:0];
  assign and_172__in0[15:0] = in_344[15:0];
  assign and_172__in1[15:0] = in_345[15:0];
  assign reg_172__in[15:0] = and_172__out[15:0];
  assign and_174__in0[15:0] = in_348[15:0];
  assign and_174__in1[15:0] = in_349[15:0];
  assign reg_174__in[15:0] = and_174__out[15:0];
  assign and_176__in0[15:0] = in_352[15:0];
  assign and_176__in1[15:0] = in_353[15:0];
  assign reg_176__in[15:0] = and_176__out[15:0];
  assign and_178__in0[15:0] = in_356[15:0];
  assign and_178__in1[15:0] = in_357[15:0];
  assign reg_178__in[15:0] = and_178__out[15:0];
  assign and_18__in0[15:0] = in_36[15:0];
  assign and_18__in1[15:0] = in_37[15:0];
  assign reg_18__in[15:0] = and_18__out[15:0];
  assign and_180__in0[15:0] = in_360[15:0];
  assign and_180__in1[15:0] = in_361[15:0];
  assign reg_180__in[15:0] = and_180__out[15:0];
  assign and_182__in0[15:0] = in_364[15:0];
  assign and_182__in1[15:0] = in_365[15:0];
  assign reg_182__in[15:0] = and_182__out[15:0];
  assign and_184__in0[15:0] = in_368[15:0];
  assign and_184__in1[15:0] = in_369[15:0];
  assign reg_184__in[15:0] = and_184__out[15:0];
  assign and_186__in0[15:0] = in_372[15:0];
  assign and_186__in1[15:0] = in_373[15:0];
  assign reg_186__in[15:0] = and_186__out[15:0];
  assign and_188__in0[15:0] = in_376[15:0];
  assign and_188__in1[15:0] = in_377[15:0];
  assign reg_188__in[15:0] = and_188__out[15:0];
  assign and_190__in0[15:0] = in_380[15:0];
  assign and_190__in1[15:0] = in_381[15:0];
  assign reg_190__in[15:0] = and_190__out[15:0];
  assign and_192__in0[15:0] = in_384[15:0];
  assign and_192__in1[15:0] = in_385[15:0];
  assign reg_192__in[15:0] = and_192__out[15:0];
  assign and_194__in0[15:0] = in_388[15:0];
  assign and_194__in1[15:0] = in_389[15:0];
  assign reg_194__in[15:0] = and_194__out[15:0];
  assign and_196__in0[15:0] = in_392[15:0];
  assign and_196__in1[15:0] = in_393[15:0];
  assign reg_196__in[15:0] = and_196__out[15:0];
  assign and_198__in0[15:0] = in_396[15:0];
  assign and_198__in1[15:0] = in_397[15:0];
  assign reg_198__in[15:0] = and_198__out[15:0];
  assign and_2__in0[15:0] = in_4[15:0];
  assign and_2__in1[15:0] = in_5[15:0];
  assign reg_2__in[15:0] = and_2__out[15:0];
  assign and_20__in0[15:0] = in_40[15:0];
  assign and_20__in1[15:0] = in_41[15:0];
  assign reg_20__in[15:0] = and_20__out[15:0];
  assign and_200__in0[15:0] = in_400[15:0];
  assign and_200__in1[15:0] = in_401[15:0];
  assign reg_200__in[15:0] = and_200__out[15:0];
  assign and_202__in0[15:0] = in_404[15:0];
  assign and_202__in1[15:0] = in_405[15:0];
  assign reg_202__in[15:0] = and_202__out[15:0];
  assign and_204__in0[15:0] = in_408[15:0];
  assign and_204__in1[15:0] = in_409[15:0];
  assign reg_204__in[15:0] = and_204__out[15:0];
  assign and_206__in0[15:0] = in_412[15:0];
  assign and_206__in1[15:0] = in_413[15:0];
  assign reg_206__in[15:0] = and_206__out[15:0];
  assign and_208__in0[15:0] = in_416[15:0];
  assign and_208__in1[15:0] = in_417[15:0];
  assign reg_208__in[15:0] = and_208__out[15:0];
  assign and_210__in0[15:0] = in_420[15:0];
  assign and_210__in1[15:0] = in_421[15:0];
  assign reg_210__in[15:0] = and_210__out[15:0];
  assign and_212__in0[15:0] = in_424[15:0];
  assign and_212__in1[15:0] = in_425[15:0];
  assign reg_212__in[15:0] = and_212__out[15:0];
  assign and_214__in0[15:0] = in_428[15:0];
  assign and_214__in1[15:0] = in_429[15:0];
  assign reg_214__in[15:0] = and_214__out[15:0];
  assign and_216__in0[15:0] = in_432[15:0];
  assign and_216__in1[15:0] = in_433[15:0];
  assign reg_216__in[15:0] = and_216__out[15:0];
  assign and_218__in0[15:0] = in_436[15:0];
  assign and_218__in1[15:0] = in_437[15:0];
  assign reg_218__in[15:0] = and_218__out[15:0];
  assign and_22__in0[15:0] = in_44[15:0];
  assign and_22__in1[15:0] = in_45[15:0];
  assign reg_22__in[15:0] = and_22__out[15:0];
  assign and_220__in0[15:0] = in_440[15:0];
  assign and_220__in1[15:0] = in_441[15:0];
  assign reg_220__in[15:0] = and_220__out[15:0];
  assign and_222__in0[15:0] = in_444[15:0];
  assign and_222__in1[15:0] = in_445[15:0];
  assign reg_222__in[15:0] = and_222__out[15:0];
  assign and_224__in0[15:0] = in_448[15:0];
  assign and_224__in1[15:0] = in_449[15:0];
  assign reg_224__in[15:0] = and_224__out[15:0];
  assign and_226__in0[15:0] = in_452[15:0];
  assign and_226__in1[15:0] = in_453[15:0];
  assign reg_226__in[15:0] = and_226__out[15:0];
  assign and_228__in0[15:0] = in_456[15:0];
  assign and_228__in1[15:0] = in_457[15:0];
  assign reg_228__in[15:0] = and_228__out[15:0];
  assign and_230__in0[15:0] = in_460[15:0];
  assign and_230__in1[15:0] = in_461[15:0];
  assign reg_230__in[15:0] = and_230__out[15:0];
  assign and_232__in0[15:0] = in_464[15:0];
  assign and_232__in1[15:0] = in_465[15:0];
  assign reg_232__in[15:0] = and_232__out[15:0];
  assign and_234__in0[15:0] = in_468[15:0];
  assign and_234__in1[15:0] = in_469[15:0];
  assign reg_234__in[15:0] = and_234__out[15:0];
  assign and_236__in0[15:0] = in_472[15:0];
  assign and_236__in1[15:0] = in_473[15:0];
  assign reg_236__in[15:0] = and_236__out[15:0];
  assign and_238__in0[15:0] = in_476[15:0];
  assign and_238__in1[15:0] = in_477[15:0];
  assign reg_238__in[15:0] = and_238__out[15:0];
  assign and_24__in0[15:0] = in_48[15:0];
  assign and_24__in1[15:0] = in_49[15:0];
  assign reg_24__in[15:0] = and_24__out[15:0];
  assign and_240__in0[15:0] = in_480[15:0];
  assign and_240__in1[15:0] = in_481[15:0];
  assign reg_240__in[15:0] = and_240__out[15:0];
  assign and_242__in0[15:0] = in_484[15:0];
  assign and_242__in1[15:0] = in_485[15:0];
  assign reg_242__in[15:0] = and_242__out[15:0];
  assign and_244__in0[15:0] = in_488[15:0];
  assign and_244__in1[15:0] = in_489[15:0];
  assign reg_244__in[15:0] = and_244__out[15:0];
  assign and_246__in0[15:0] = in_492[15:0];
  assign and_246__in1[15:0] = in_493[15:0];
  assign reg_246__in[15:0] = and_246__out[15:0];
  assign and_248__in0[15:0] = in_496[15:0];
  assign and_248__in1[15:0] = in_497[15:0];
  assign reg_248__in[15:0] = and_248__out[15:0];
  assign and_250__in0[15:0] = in_500[15:0];
  assign and_250__in1[15:0] = in_501[15:0];
  assign reg_250__in[15:0] = and_250__out[15:0];
  assign and_252__in0[15:0] = in_504[15:0];
  assign and_252__in1[15:0] = in_505[15:0];
  assign reg_252__in[15:0] = and_252__out[15:0];
  assign and_254__in0[15:0] = in_508[15:0];
  assign and_254__in1[15:0] = in_509[15:0];
  assign reg_254__in[15:0] = and_254__out[15:0];
  assign and_256__in0[15:0] = in_512[15:0];
  assign and_256__in1[15:0] = in_513[15:0];
  assign reg_256__in[15:0] = and_256__out[15:0];
  assign and_258__in0[15:0] = in_516[15:0];
  assign and_258__in1[15:0] = in_517[15:0];
  assign reg_258__in[15:0] = and_258__out[15:0];
  assign and_26__in0[15:0] = in_52[15:0];
  assign and_26__in1[15:0] = in_53[15:0];
  assign reg_26__in[15:0] = and_26__out[15:0];
  assign and_260__in0[15:0] = in_520[15:0];
  assign and_260__in1[15:0] = in_521[15:0];
  assign reg_260__in[15:0] = and_260__out[15:0];
  assign and_262__in0[15:0] = in_524[15:0];
  assign and_262__in1[15:0] = in_525[15:0];
  assign reg_262__in[15:0] = and_262__out[15:0];
  assign and_264__in0[15:0] = in_528[15:0];
  assign and_264__in1[15:0] = in_529[15:0];
  assign reg_264__in[15:0] = and_264__out[15:0];
  assign and_266__in0[15:0] = in_532[15:0];
  assign and_266__in1[15:0] = in_533[15:0];
  assign reg_266__in[15:0] = and_266__out[15:0];
  assign and_268__in0[15:0] = in_536[15:0];
  assign and_268__in1[15:0] = in_537[15:0];
  assign reg_268__in[15:0] = and_268__out[15:0];
  assign and_270__in0[15:0] = in_540[15:0];
  assign and_270__in1[15:0] = in_541[15:0];
  assign reg_270__in[15:0] = and_270__out[15:0];
  assign and_272__in0[15:0] = in_544[15:0];
  assign and_272__in1[15:0] = in_545[15:0];
  assign reg_272__in[15:0] = and_272__out[15:0];
  assign and_274__in0[15:0] = in_548[15:0];
  assign and_274__in1[15:0] = in_549[15:0];
  assign reg_274__in[15:0] = and_274__out[15:0];
  assign and_276__in0[15:0] = in_552[15:0];
  assign and_276__in1[15:0] = in_553[15:0];
  assign reg_276__in[15:0] = and_276__out[15:0];
  assign and_278__in0[15:0] = in_556[15:0];
  assign and_278__in1[15:0] = in_557[15:0];
  assign reg_278__in[15:0] = and_278__out[15:0];
  assign and_28__in0[15:0] = in_56[15:0];
  assign and_28__in1[15:0] = in_57[15:0];
  assign reg_28__in[15:0] = and_28__out[15:0];
  assign and_280__in0[15:0] = in_560[15:0];
  assign and_280__in1[15:0] = in_561[15:0];
  assign reg_280__in[15:0] = and_280__out[15:0];
  assign and_282__in0[15:0] = in_564[15:0];
  assign and_282__in1[15:0] = in_565[15:0];
  assign reg_282__in[15:0] = and_282__out[15:0];
  assign and_284__in0[15:0] = in_568[15:0];
  assign and_284__in1[15:0] = in_569[15:0];
  assign reg_284__in[15:0] = and_284__out[15:0];
  assign and_286__in0[15:0] = in_572[15:0];
  assign and_286__in1[15:0] = in_573[15:0];
  assign reg_286__in[15:0] = and_286__out[15:0];
  assign and_288__in0[15:0] = in_576[15:0];
  assign and_288__in1[15:0] = in_577[15:0];
  assign reg_288__in[15:0] = and_288__out[15:0];
  assign and_290__in0[15:0] = in_580[15:0];
  assign and_290__in1[15:0] = in_581[15:0];
  assign reg_290__in[15:0] = and_290__out[15:0];
  assign and_292__in0[15:0] = in_584[15:0];
  assign and_292__in1[15:0] = in_585[15:0];
  assign reg_292__in[15:0] = and_292__out[15:0];
  assign and_294__in0[15:0] = in_588[15:0];
  assign and_294__in1[15:0] = in_589[15:0];
  assign reg_294__in[15:0] = and_294__out[15:0];
  assign and_296__in0[15:0] = in_592[15:0];
  assign and_296__in1[15:0] = in_593[15:0];
  assign reg_296__in[15:0] = and_296__out[15:0];
  assign and_298__in0[15:0] = in_596[15:0];
  assign and_298__in1[15:0] = in_597[15:0];
  assign reg_298__in[15:0] = and_298__out[15:0];
  assign and_30__in0[15:0] = in_60[15:0];
  assign and_30__in1[15:0] = in_61[15:0];
  assign reg_30__in[15:0] = and_30__out[15:0];
  assign and_300__in0[15:0] = in_600[15:0];
  assign and_300__in1[15:0] = in_601[15:0];
  assign reg_300__in[15:0] = and_300__out[15:0];
  assign and_302__in0[15:0] = in_604[15:0];
  assign and_302__in1[15:0] = in_605[15:0];
  assign reg_302__in[15:0] = and_302__out[15:0];
  assign and_304__in0[15:0] = in_608[15:0];
  assign and_304__in1[15:0] = in_609[15:0];
  assign reg_304__in[15:0] = and_304__out[15:0];
  assign and_306__in0[15:0] = in_612[15:0];
  assign and_306__in1[15:0] = in_613[15:0];
  assign reg_306__in[15:0] = and_306__out[15:0];
  assign and_308__in0[15:0] = in_616[15:0];
  assign and_308__in1[15:0] = in_617[15:0];
  assign reg_308__in[15:0] = and_308__out[15:0];
  assign and_310__in0[15:0] = in_620[15:0];
  assign and_310__in1[15:0] = in_621[15:0];
  assign reg_310__in[15:0] = and_310__out[15:0];
  assign and_312__in0[15:0] = in_624[15:0];
  assign and_312__in1[15:0] = in_625[15:0];
  assign reg_312__in[15:0] = and_312__out[15:0];
  assign and_314__in0[15:0] = in_628[15:0];
  assign and_314__in1[15:0] = in_629[15:0];
  assign reg_314__in[15:0] = and_314__out[15:0];
  assign and_316__in0[15:0] = in_632[15:0];
  assign and_316__in1[15:0] = in_633[15:0];
  assign reg_316__in[15:0] = and_316__out[15:0];
  assign and_318__in0[15:0] = in_636[15:0];
  assign and_318__in1[15:0] = in_637[15:0];
  assign reg_318__in[15:0] = and_318__out[15:0];
  assign and_32__in0[15:0] = in_64[15:0];
  assign and_32__in1[15:0] = in_65[15:0];
  assign reg_32__in[15:0] = and_32__out[15:0];
  assign and_320__in0[15:0] = in_640[15:0];
  assign and_320__in1[15:0] = in_641[15:0];
  assign reg_320__in[15:0] = and_320__out[15:0];
  assign and_322__in0[15:0] = in_644[15:0];
  assign and_322__in1[15:0] = in_645[15:0];
  assign reg_322__in[15:0] = and_322__out[15:0];
  assign and_324__in0[15:0] = in_648[15:0];
  assign and_324__in1[15:0] = in_649[15:0];
  assign reg_324__in[15:0] = and_324__out[15:0];
  assign and_326__in0[15:0] = in_652[15:0];
  assign and_326__in1[15:0] = in_653[15:0];
  assign reg_326__in[15:0] = and_326__out[15:0];
  assign and_328__in0[15:0] = in_656[15:0];
  assign and_328__in1[15:0] = in_657[15:0];
  assign reg_328__in[15:0] = and_328__out[15:0];
  assign and_330__in0[15:0] = in_660[15:0];
  assign and_330__in1[15:0] = in_661[15:0];
  assign reg_330__in[15:0] = and_330__out[15:0];
  assign and_332__in0[15:0] = in_664[15:0];
  assign and_332__in1[15:0] = in_665[15:0];
  assign reg_332__in[15:0] = and_332__out[15:0];
  assign and_334__in0[15:0] = in_668[15:0];
  assign and_334__in1[15:0] = in_669[15:0];
  assign reg_334__in[15:0] = and_334__out[15:0];
  assign and_336__in0[15:0] = in_672[15:0];
  assign and_336__in1[15:0] = in_673[15:0];
  assign reg_336__in[15:0] = and_336__out[15:0];
  assign and_338__in0[15:0] = in_676[15:0];
  assign and_338__in1[15:0] = in_677[15:0];
  assign reg_338__in[15:0] = and_338__out[15:0];
  assign and_34__in0[15:0] = in_68[15:0];
  assign and_34__in1[15:0] = in_69[15:0];
  assign reg_34__in[15:0] = and_34__out[15:0];
  assign and_340__in0[15:0] = in_680[15:0];
  assign and_340__in1[15:0] = in_681[15:0];
  assign reg_340__in[15:0] = and_340__out[15:0];
  assign and_342__in0[15:0] = in_684[15:0];
  assign and_342__in1[15:0] = in_685[15:0];
  assign reg_342__in[15:0] = and_342__out[15:0];
  assign and_344__in0[15:0] = in_688[15:0];
  assign and_344__in1[15:0] = in_689[15:0];
  assign reg_344__in[15:0] = and_344__out[15:0];
  assign and_346__in0[15:0] = in_692[15:0];
  assign and_346__in1[15:0] = in_693[15:0];
  assign reg_346__in[15:0] = and_346__out[15:0];
  assign and_348__in0[15:0] = in_696[15:0];
  assign and_348__in1[15:0] = in_697[15:0];
  assign reg_348__in[15:0] = and_348__out[15:0];
  assign and_350__in0[15:0] = in_700[15:0];
  assign and_350__in1[15:0] = in_701[15:0];
  assign reg_350__in[15:0] = and_350__out[15:0];
  assign and_352__in0[15:0] = in_704[15:0];
  assign and_352__in1[15:0] = in_705[15:0];
  assign reg_352__in[15:0] = and_352__out[15:0];
  assign and_354__in0[15:0] = in_708[15:0];
  assign and_354__in1[15:0] = in_709[15:0];
  assign reg_354__in[15:0] = and_354__out[15:0];
  assign and_356__in0[15:0] = in_712[15:0];
  assign and_356__in1[15:0] = in_713[15:0];
  assign reg_356__in[15:0] = and_356__out[15:0];
  assign and_358__in0[15:0] = in_716[15:0];
  assign and_358__in1[15:0] = in_717[15:0];
  assign reg_358__in[15:0] = and_358__out[15:0];
  assign and_36__in0[15:0] = in_72[15:0];
  assign and_36__in1[15:0] = in_73[15:0];
  assign reg_36__in[15:0] = and_36__out[15:0];
  assign and_360__in0[15:0] = in_720[15:0];
  assign and_360__in1[15:0] = in_721[15:0];
  assign reg_360__in[15:0] = and_360__out[15:0];
  assign and_362__in0[15:0] = in_724[15:0];
  assign and_362__in1[15:0] = in_725[15:0];
  assign reg_362__in[15:0] = and_362__out[15:0];
  assign and_364__in0[15:0] = in_728[15:0];
  assign and_364__in1[15:0] = in_729[15:0];
  assign reg_364__in[15:0] = and_364__out[15:0];
  assign and_366__in0[15:0] = in_732[15:0];
  assign and_366__in1[15:0] = in_733[15:0];
  assign reg_366__in[15:0] = and_366__out[15:0];
  assign and_368__in0[15:0] = in_736[15:0];
  assign and_368__in1[15:0] = in_737[15:0];
  assign reg_368__in[15:0] = and_368__out[15:0];
  assign and_370__in0[15:0] = in_740[15:0];
  assign and_370__in1[15:0] = in_741[15:0];
  assign reg_370__in[15:0] = and_370__out[15:0];
  assign and_372__in0[15:0] = in_744[15:0];
  assign and_372__in1[15:0] = in_745[15:0];
  assign reg_372__in[15:0] = and_372__out[15:0];
  assign and_374__in0[15:0] = in_748[15:0];
  assign and_374__in1[15:0] = in_749[15:0];
  assign reg_374__in[15:0] = and_374__out[15:0];
  assign and_376__in0[15:0] = in_752[15:0];
  assign and_376__in1[15:0] = in_753[15:0];
  assign reg_376__in[15:0] = and_376__out[15:0];
  assign and_378__in0[15:0] = in_756[15:0];
  assign and_378__in1[15:0] = in_757[15:0];
  assign reg_378__in[15:0] = and_378__out[15:0];
  assign and_38__in0[15:0] = in_76[15:0];
  assign and_38__in1[15:0] = in_77[15:0];
  assign reg_38__in[15:0] = and_38__out[15:0];
  assign and_380__in0[15:0] = in_760[15:0];
  assign and_380__in1[15:0] = in_761[15:0];
  assign reg_380__in[15:0] = and_380__out[15:0];
  assign and_382__in0[15:0] = in_764[15:0];
  assign and_382__in1[15:0] = in_765[15:0];
  assign reg_382__in[15:0] = and_382__out[15:0];
  assign and_384__in0[15:0] = in_768[15:0];
  assign and_384__in1[15:0] = in_769[15:0];
  assign reg_384__in[15:0] = and_384__out[15:0];
  assign and_386__in0[15:0] = in_772[15:0];
  assign and_386__in1[15:0] = in_773[15:0];
  assign reg_386__in[15:0] = and_386__out[15:0];
  assign and_388__in0[15:0] = in_776[15:0];
  assign and_388__in1[15:0] = in_777[15:0];
  assign reg_388__in[15:0] = and_388__out[15:0];
  assign and_390__in0[15:0] = in_780[15:0];
  assign and_390__in1[15:0] = in_781[15:0];
  assign reg_390__in[15:0] = and_390__out[15:0];
  assign and_392__in0[15:0] = in_784[15:0];
  assign and_392__in1[15:0] = in_785[15:0];
  assign reg_392__in[15:0] = and_392__out[15:0];
  assign and_394__in0[15:0] = in_788[15:0];
  assign and_394__in1[15:0] = in_789[15:0];
  assign reg_394__in[15:0] = and_394__out[15:0];
  assign and_396__in0[15:0] = in_792[15:0];
  assign and_396__in1[15:0] = in_793[15:0];
  assign reg_396__in[15:0] = and_396__out[15:0];
  assign and_398__in0[15:0] = in_796[15:0];
  assign and_398__in1[15:0] = in_797[15:0];
  assign reg_398__in[15:0] = and_398__out[15:0];
  assign and_4__in0[15:0] = in_8[15:0];
  assign and_4__in1[15:0] = in_9[15:0];
  assign reg_4__in[15:0] = and_4__out[15:0];
  assign and_40__in0[15:0] = in_80[15:0];
  assign and_40__in1[15:0] = in_81[15:0];
  assign reg_40__in[15:0] = and_40__out[15:0];
  assign and_400__in0[15:0] = in_800[15:0];
  assign and_400__in1[15:0] = in_801[15:0];
  assign reg_400__in[15:0] = and_400__out[15:0];
  assign and_402__in0[15:0] = in_804[15:0];
  assign and_402__in1[15:0] = in_805[15:0];
  assign reg_402__in[15:0] = and_402__out[15:0];
  assign and_404__in0[15:0] = in_808[15:0];
  assign and_404__in1[15:0] = in_809[15:0];
  assign reg_404__in[15:0] = and_404__out[15:0];
  assign and_406__in0[15:0] = in_812[15:0];
  assign and_406__in1[15:0] = in_813[15:0];
  assign reg_406__in[15:0] = and_406__out[15:0];
  assign and_408__in0[15:0] = in_816[15:0];
  assign and_408__in1[15:0] = in_817[15:0];
  assign reg_408__in[15:0] = and_408__out[15:0];
  assign and_410__in0[15:0] = in_820[15:0];
  assign and_410__in1[15:0] = in_821[15:0];
  assign reg_410__in[15:0] = and_410__out[15:0];
  assign and_412__in0[15:0] = in_824[15:0];
  assign and_412__in1[15:0] = in_825[15:0];
  assign reg_412__in[15:0] = and_412__out[15:0];
  assign and_414__in0[15:0] = in_828[15:0];
  assign and_414__in1[15:0] = in_829[15:0];
  assign reg_414__in[15:0] = and_414__out[15:0];
  assign and_416__in0[15:0] = in_832[15:0];
  assign and_416__in1[15:0] = in_833[15:0];
  assign reg_416__in[15:0] = and_416__out[15:0];
  assign and_418__in0[15:0] = in_836[15:0];
  assign and_418__in1[15:0] = in_837[15:0];
  assign reg_418__in[15:0] = and_418__out[15:0];
  assign and_42__in0[15:0] = in_84[15:0];
  assign and_42__in1[15:0] = in_85[15:0];
  assign reg_42__in[15:0] = and_42__out[15:0];
  assign and_420__in0[15:0] = in_840[15:0];
  assign and_420__in1[15:0] = in_841[15:0];
  assign reg_420__in[15:0] = and_420__out[15:0];
  assign and_422__in0[15:0] = in_844[15:0];
  assign and_422__in1[15:0] = in_845[15:0];
  assign reg_422__in[15:0] = and_422__out[15:0];
  assign and_424__in0[15:0] = in_848[15:0];
  assign and_424__in1[15:0] = in_849[15:0];
  assign reg_424__in[15:0] = and_424__out[15:0];
  assign and_426__in0[15:0] = in_852[15:0];
  assign and_426__in1[15:0] = in_853[15:0];
  assign reg_426__in[15:0] = and_426__out[15:0];
  assign and_428__in0[15:0] = in_856[15:0];
  assign and_428__in1[15:0] = in_857[15:0];
  assign reg_428__in[15:0] = and_428__out[15:0];
  assign and_430__in0[15:0] = in_860[15:0];
  assign and_430__in1[15:0] = in_861[15:0];
  assign reg_430__in[15:0] = and_430__out[15:0];
  assign and_432__in0[15:0] = in_864[15:0];
  assign and_432__in1[15:0] = in_865[15:0];
  assign reg_432__in[15:0] = and_432__out[15:0];
  assign and_434__in0[15:0] = in_868[15:0];
  assign and_434__in1[15:0] = in_869[15:0];
  assign reg_434__in[15:0] = and_434__out[15:0];
  assign and_436__in0[15:0] = in_872[15:0];
  assign and_436__in1[15:0] = in_873[15:0];
  assign reg_436__in[15:0] = and_436__out[15:0];
  assign and_438__in0[15:0] = in_876[15:0];
  assign and_438__in1[15:0] = in_877[15:0];
  assign reg_438__in[15:0] = and_438__out[15:0];
  assign and_44__in0[15:0] = in_88[15:0];
  assign and_44__in1[15:0] = in_89[15:0];
  assign reg_44__in[15:0] = and_44__out[15:0];
  assign and_440__in0[15:0] = in_880[15:0];
  assign and_440__in1[15:0] = in_881[15:0];
  assign reg_440__in[15:0] = and_440__out[15:0];
  assign and_442__in0[15:0] = in_884[15:0];
  assign and_442__in1[15:0] = in_885[15:0];
  assign reg_442__in[15:0] = and_442__out[15:0];
  assign and_444__in0[15:0] = in_888[15:0];
  assign and_444__in1[15:0] = in_889[15:0];
  assign reg_444__in[15:0] = and_444__out[15:0];
  assign and_446__in0[15:0] = in_892[15:0];
  assign and_446__in1[15:0] = in_893[15:0];
  assign reg_446__in[15:0] = and_446__out[15:0];
  assign and_448__in0[15:0] = in_896[15:0];
  assign and_448__in1[15:0] = in_897[15:0];
  assign reg_448__in[15:0] = and_448__out[15:0];
  assign and_450__in0[15:0] = in_900[15:0];
  assign and_450__in1[15:0] = in_901[15:0];
  assign reg_450__in[15:0] = and_450__out[15:0];
  assign and_452__in0[15:0] = in_904[15:0];
  assign and_452__in1[15:0] = in_905[15:0];
  assign reg_452__in[15:0] = and_452__out[15:0];
  assign and_454__in0[15:0] = in_908[15:0];
  assign and_454__in1[15:0] = in_909[15:0];
  assign reg_454__in[15:0] = and_454__out[15:0];
  assign and_456__in0[15:0] = in_912[15:0];
  assign and_456__in1[15:0] = in_913[15:0];
  assign reg_456__in[15:0] = and_456__out[15:0];
  assign and_458__in0[15:0] = in_916[15:0];
  assign and_458__in1[15:0] = in_917[15:0];
  assign reg_458__in[15:0] = and_458__out[15:0];
  assign and_46__in0[15:0] = in_92[15:0];
  assign and_46__in1[15:0] = in_93[15:0];
  assign reg_46__in[15:0] = and_46__out[15:0];
  assign and_460__in0[15:0] = in_920[15:0];
  assign and_460__in1[15:0] = in_921[15:0];
  assign reg_460__in[15:0] = and_460__out[15:0];
  assign and_462__in0[15:0] = in_924[15:0];
  assign and_462__in1[15:0] = in_925[15:0];
  assign reg_462__in[15:0] = and_462__out[15:0];
  assign and_464__in0[15:0] = in_928[15:0];
  assign and_464__in1[15:0] = in_929[15:0];
  assign reg_464__in[15:0] = and_464__out[15:0];
  assign and_466__in0[15:0] = in_932[15:0];
  assign and_466__in1[15:0] = in_933[15:0];
  assign reg_466__in[15:0] = and_466__out[15:0];
  assign and_468__in0[15:0] = in_936[15:0];
  assign and_468__in1[15:0] = in_937[15:0];
  assign reg_468__in[15:0] = and_468__out[15:0];
  assign and_470__in0[15:0] = in_940[15:0];
  assign and_470__in1[15:0] = in_941[15:0];
  assign reg_470__in[15:0] = and_470__out[15:0];
  assign and_472__in0[15:0] = in_944[15:0];
  assign and_472__in1[15:0] = in_945[15:0];
  assign reg_472__in[15:0] = and_472__out[15:0];
  assign and_474__in0[15:0] = in_948[15:0];
  assign and_474__in1[15:0] = in_949[15:0];
  assign reg_474__in[15:0] = and_474__out[15:0];
  assign and_476__in0[15:0] = in_952[15:0];
  assign and_476__in1[15:0] = in_953[15:0];
  assign reg_476__in[15:0] = and_476__out[15:0];
  assign and_478__in0[15:0] = in_956[15:0];
  assign and_478__in1[15:0] = in_957[15:0];
  assign reg_478__in[15:0] = and_478__out[15:0];
  assign and_48__in0[15:0] = in_96[15:0];
  assign and_48__in1[15:0] = in_97[15:0];
  assign reg_48__in[15:0] = and_48__out[15:0];
  assign and_480__in0[15:0] = in_960[15:0];
  assign and_480__in1[15:0] = in_961[15:0];
  assign reg_480__in[15:0] = and_480__out[15:0];
  assign and_482__in0[15:0] = in_964[15:0];
  assign and_482__in1[15:0] = in_965[15:0];
  assign reg_482__in[15:0] = and_482__out[15:0];
  assign and_484__in0[15:0] = in_968[15:0];
  assign and_484__in1[15:0] = in_969[15:0];
  assign reg_484__in[15:0] = and_484__out[15:0];
  assign and_486__in0[15:0] = in_972[15:0];
  assign and_486__in1[15:0] = in_973[15:0];
  assign reg_486__in[15:0] = and_486__out[15:0];
  assign and_488__in0[15:0] = in_976[15:0];
  assign and_488__in1[15:0] = in_977[15:0];
  assign reg_488__in[15:0] = and_488__out[15:0];
  assign and_490__in0[15:0] = in_980[15:0];
  assign and_490__in1[15:0] = in_981[15:0];
  assign reg_490__in[15:0] = and_490__out[15:0];
  assign and_492__in0[15:0] = in_984[15:0];
  assign and_492__in1[15:0] = in_985[15:0];
  assign reg_492__in[15:0] = and_492__out[15:0];
  assign and_494__in0[15:0] = in_988[15:0];
  assign and_494__in1[15:0] = in_989[15:0];
  assign reg_494__in[15:0] = and_494__out[15:0];
  assign and_496__in0[15:0] = in_992[15:0];
  assign and_496__in1[15:0] = in_993[15:0];
  assign reg_496__in[15:0] = and_496__out[15:0];
  assign and_498__in0[15:0] = in_996[15:0];
  assign and_498__in1[15:0] = in_997[15:0];
  assign reg_498__in[15:0] = and_498__out[15:0];
  assign and_50__in0[15:0] = in_100[15:0];
  assign and_50__in1[15:0] = in_101[15:0];
  assign reg_50__in[15:0] = and_50__out[15:0];
  assign and_500__in0[15:0] = in_1000[15:0];
  assign and_500__in1[15:0] = in_1001[15:0];
  assign reg_500__in[15:0] = and_500__out[15:0];
  assign and_502__in0[15:0] = in_1004[15:0];
  assign and_502__in1[15:0] = in_1005[15:0];
  assign reg_502__in[15:0] = and_502__out[15:0];
  assign and_504__in0[15:0] = in_1008[15:0];
  assign and_504__in1[15:0] = in_1009[15:0];
  assign reg_504__in[15:0] = and_504__out[15:0];
  assign and_506__in0[15:0] = in_1012[15:0];
  assign and_506__in1[15:0] = in_1013[15:0];
  assign reg_506__in[15:0] = and_506__out[15:0];
  assign and_508__in0[15:0] = in_1016[15:0];
  assign and_508__in1[15:0] = in_1017[15:0];
  assign reg_508__in[15:0] = and_508__out[15:0];
  assign and_510__in0[15:0] = in_1020[15:0];
  assign and_510__in1[15:0] = in_1021[15:0];
  assign reg_510__in[15:0] = and_510__out[15:0];
  assign and_512__in0[15:0] = in_1024[15:0];
  assign and_512__in1[15:0] = in_1025[15:0];
  assign reg_512__in[15:0] = and_512__out[15:0];
  assign and_514__in0[15:0] = in_1028[15:0];
  assign and_514__in1[15:0] = in_1029[15:0];
  assign reg_514__in[15:0] = and_514__out[15:0];
  assign and_516__in0[15:0] = in_1032[15:0];
  assign and_516__in1[15:0] = in_1033[15:0];
  assign reg_516__in[15:0] = and_516__out[15:0];
  assign and_518__in0[15:0] = in_1036[15:0];
  assign and_518__in1[15:0] = in_1037[15:0];
  assign reg_518__in[15:0] = and_518__out[15:0];
  assign and_52__in0[15:0] = in_104[15:0];
  assign and_52__in1[15:0] = in_105[15:0];
  assign reg_52__in[15:0] = and_52__out[15:0];
  assign and_520__in0[15:0] = in_1040[15:0];
  assign and_520__in1[15:0] = in_1041[15:0];
  assign reg_520__in[15:0] = and_520__out[15:0];
  assign and_522__in0[15:0] = in_1044[15:0];
  assign and_522__in1[15:0] = in_1045[15:0];
  assign reg_522__in[15:0] = and_522__out[15:0];
  assign and_524__in0[15:0] = in_1048[15:0];
  assign and_524__in1[15:0] = in_1049[15:0];
  assign reg_524__in[15:0] = and_524__out[15:0];
  assign and_526__in0[15:0] = in_1052[15:0];
  assign and_526__in1[15:0] = in_1053[15:0];
  assign reg_526__in[15:0] = and_526__out[15:0];
  assign and_528__in0[15:0] = in_1056[15:0];
  assign and_528__in1[15:0] = in_1057[15:0];
  assign reg_528__in[15:0] = and_528__out[15:0];
  assign and_530__in0[15:0] = in_1060[15:0];
  assign and_530__in1[15:0] = in_1061[15:0];
  assign reg_530__in[15:0] = and_530__out[15:0];
  assign and_532__in0[15:0] = in_1064[15:0];
  assign and_532__in1[15:0] = in_1065[15:0];
  assign reg_532__in[15:0] = and_532__out[15:0];
  assign and_534__in0[15:0] = in_1068[15:0];
  assign and_534__in1[15:0] = in_1069[15:0];
  assign reg_534__in[15:0] = and_534__out[15:0];
  assign and_536__in0[15:0] = in_1072[15:0];
  assign and_536__in1[15:0] = in_1073[15:0];
  assign reg_536__in[15:0] = and_536__out[15:0];
  assign and_538__in0[15:0] = in_1076[15:0];
  assign and_538__in1[15:0] = in_1077[15:0];
  assign reg_538__in[15:0] = and_538__out[15:0];
  assign and_54__in0[15:0] = in_108[15:0];
  assign and_54__in1[15:0] = in_109[15:0];
  assign reg_54__in[15:0] = and_54__out[15:0];
  assign and_540__in0[15:0] = in_1080[15:0];
  assign and_540__in1[15:0] = in_1081[15:0];
  assign reg_540__in[15:0] = and_540__out[15:0];
  assign and_542__in0[15:0] = in_1084[15:0];
  assign and_542__in1[15:0] = in_1085[15:0];
  assign reg_542__in[15:0] = and_542__out[15:0];
  assign and_544__in0[15:0] = in_1088[15:0];
  assign and_544__in1[15:0] = in_1089[15:0];
  assign reg_544__in[15:0] = and_544__out[15:0];
  assign and_546__in0[15:0] = in_1092[15:0];
  assign and_546__in1[15:0] = in_1093[15:0];
  assign reg_546__in[15:0] = and_546__out[15:0];
  assign and_548__in0[15:0] = in_1096[15:0];
  assign and_548__in1[15:0] = in_1097[15:0];
  assign reg_548__in[15:0] = and_548__out[15:0];
  assign and_550__in0[15:0] = in_1100[15:0];
  assign and_550__in1[15:0] = in_1101[15:0];
  assign reg_550__in[15:0] = and_550__out[15:0];
  assign and_552__in0[15:0] = in_1104[15:0];
  assign and_552__in1[15:0] = in_1105[15:0];
  assign reg_552__in[15:0] = and_552__out[15:0];
  assign and_554__in0[15:0] = in_1108[15:0];
  assign and_554__in1[15:0] = in_1109[15:0];
  assign reg_554__in[15:0] = and_554__out[15:0];
  assign and_556__in0[15:0] = in_1112[15:0];
  assign and_556__in1[15:0] = in_1113[15:0];
  assign reg_556__in[15:0] = and_556__out[15:0];
  assign and_558__in0[15:0] = in_1116[15:0];
  assign and_558__in1[15:0] = in_1117[15:0];
  assign reg_558__in[15:0] = and_558__out[15:0];
  assign and_56__in0[15:0] = in_112[15:0];
  assign and_56__in1[15:0] = in_113[15:0];
  assign reg_56__in[15:0] = and_56__out[15:0];
  assign and_560__in0[15:0] = in_1120[15:0];
  assign and_560__in1[15:0] = in_1121[15:0];
  assign reg_560__in[15:0] = and_560__out[15:0];
  assign and_562__in0[15:0] = in_1124[15:0];
  assign and_562__in1[15:0] = in_1125[15:0];
  assign reg_562__in[15:0] = and_562__out[15:0];
  assign and_564__in0[15:0] = in_1128[15:0];
  assign and_564__in1[15:0] = in_1129[15:0];
  assign reg_564__in[15:0] = and_564__out[15:0];
  assign and_566__in0[15:0] = in_1132[15:0];
  assign and_566__in1[15:0] = in_1133[15:0];
  assign reg_566__in[15:0] = and_566__out[15:0];
  assign and_568__in0[15:0] = in_1136[15:0];
  assign and_568__in1[15:0] = in_1137[15:0];
  assign reg_568__in[15:0] = and_568__out[15:0];
  assign and_570__in0[15:0] = in_1140[15:0];
  assign and_570__in1[15:0] = in_1141[15:0];
  assign reg_570__in[15:0] = and_570__out[15:0];
  assign and_572__in0[15:0] = in_1144[15:0];
  assign and_572__in1[15:0] = in_1145[15:0];
  assign reg_572__in[15:0] = and_572__out[15:0];
  assign and_574__in0[15:0] = in_1148[15:0];
  assign and_574__in1[15:0] = in_1149[15:0];
  assign reg_574__in[15:0] = and_574__out[15:0];
  assign and_576__in0[15:0] = in_1152[15:0];
  assign and_576__in1[15:0] = in_1153[15:0];
  assign reg_576__in[15:0] = and_576__out[15:0];
  assign and_578__in0[15:0] = in_1156[15:0];
  assign and_578__in1[15:0] = in_1157[15:0];
  assign reg_578__in[15:0] = and_578__out[15:0];
  assign and_58__in0[15:0] = in_116[15:0];
  assign and_58__in1[15:0] = in_117[15:0];
  assign reg_58__in[15:0] = and_58__out[15:0];
  assign and_580__in0[15:0] = in_1160[15:0];
  assign and_580__in1[15:0] = in_1161[15:0];
  assign reg_580__in[15:0] = and_580__out[15:0];
  assign and_582__in0[15:0] = in_1164[15:0];
  assign and_582__in1[15:0] = in_1165[15:0];
  assign reg_582__in[15:0] = and_582__out[15:0];
  assign and_584__in0[15:0] = in_1168[15:0];
  assign and_584__in1[15:0] = in_1169[15:0];
  assign reg_584__in[15:0] = and_584__out[15:0];
  assign and_586__in0[15:0] = in_1172[15:0];
  assign and_586__in1[15:0] = in_1173[15:0];
  assign reg_586__in[15:0] = and_586__out[15:0];
  assign and_588__in0[15:0] = in_1176[15:0];
  assign and_588__in1[15:0] = in_1177[15:0];
  assign reg_588__in[15:0] = and_588__out[15:0];
  assign and_590__in0[15:0] = in_1180[15:0];
  assign and_590__in1[15:0] = in_1181[15:0];
  assign reg_590__in[15:0] = and_590__out[15:0];
  assign and_592__in0[15:0] = in_1184[15:0];
  assign and_592__in1[15:0] = in_1185[15:0];
  assign reg_592__in[15:0] = and_592__out[15:0];
  assign and_594__in0[15:0] = in_1188[15:0];
  assign and_594__in1[15:0] = in_1189[15:0];
  assign reg_594__in[15:0] = and_594__out[15:0];
  assign and_596__in0[15:0] = in_1192[15:0];
  assign and_596__in1[15:0] = in_1193[15:0];
  assign reg_596__in[15:0] = and_596__out[15:0];
  assign and_598__in0[15:0] = in_1196[15:0];
  assign and_598__in1[15:0] = in_1197[15:0];
  assign reg_598__in[15:0] = and_598__out[15:0];
  assign and_6__in0[15:0] = in_12[15:0];
  assign and_6__in1[15:0] = in_13[15:0];
  assign reg_6__in[15:0] = and_6__out[15:0];
  assign and_60__in0[15:0] = in_120[15:0];
  assign and_60__in1[15:0] = in_121[15:0];
  assign reg_60__in[15:0] = and_60__out[15:0];
  assign and_600__in0[15:0] = in_1200[15:0];
  assign and_600__in1[15:0] = in_1201[15:0];
  assign reg_600__in[15:0] = and_600__out[15:0];
  assign and_602__in0[15:0] = in_1204[15:0];
  assign and_602__in1[15:0] = in_1205[15:0];
  assign reg_602__in[15:0] = and_602__out[15:0];
  assign and_604__in0[15:0] = in_1208[15:0];
  assign and_604__in1[15:0] = in_1209[15:0];
  assign reg_604__in[15:0] = and_604__out[15:0];
  assign and_606__in0[15:0] = in_1212[15:0];
  assign and_606__in1[15:0] = in_1213[15:0];
  assign reg_606__in[15:0] = and_606__out[15:0];
  assign and_608__in0[15:0] = in_1216[15:0];
  assign and_608__in1[15:0] = in_1217[15:0];
  assign reg_608__in[15:0] = and_608__out[15:0];
  assign and_610__in0[15:0] = in_1220[15:0];
  assign and_610__in1[15:0] = in_1221[15:0];
  assign reg_610__in[15:0] = and_610__out[15:0];
  assign and_612__in0[15:0] = in_1224[15:0];
  assign and_612__in1[15:0] = in_1225[15:0];
  assign reg_612__in[15:0] = and_612__out[15:0];
  assign and_614__in0[15:0] = in_1228[15:0];
  assign and_614__in1[15:0] = in_1229[15:0];
  assign reg_614__in[15:0] = and_614__out[15:0];
  assign and_616__in0[15:0] = in_1232[15:0];
  assign and_616__in1[15:0] = in_1233[15:0];
  assign reg_616__in[15:0] = and_616__out[15:0];
  assign and_618__in0[15:0] = in_1236[15:0];
  assign and_618__in1[15:0] = in_1237[15:0];
  assign reg_618__in[15:0] = and_618__out[15:0];
  assign and_62__in0[15:0] = in_124[15:0];
  assign and_62__in1[15:0] = in_125[15:0];
  assign reg_62__in[15:0] = and_62__out[15:0];
  assign and_620__in0[15:0] = in_1240[15:0];
  assign and_620__in1[15:0] = in_1241[15:0];
  assign reg_620__in[15:0] = and_620__out[15:0];
  assign and_622__in0[15:0] = in_1244[15:0];
  assign and_622__in1[15:0] = in_1245[15:0];
  assign reg_622__in[15:0] = and_622__out[15:0];
  assign and_624__in0[15:0] = in_1248[15:0];
  assign and_624__in1[15:0] = in_1249[15:0];
  assign reg_624__in[15:0] = and_624__out[15:0];
  assign and_626__in0[15:0] = in_1252[15:0];
  assign and_626__in1[15:0] = in_1253[15:0];
  assign reg_626__in[15:0] = and_626__out[15:0];
  assign and_628__in0[15:0] = in_1256[15:0];
  assign and_628__in1[15:0] = in_1257[15:0];
  assign reg_628__in[15:0] = and_628__out[15:0];
  assign and_630__in0[15:0] = in_1260[15:0];
  assign and_630__in1[15:0] = in_1261[15:0];
  assign reg_630__in[15:0] = and_630__out[15:0];
  assign and_632__in0[15:0] = in_1264[15:0];
  assign and_632__in1[15:0] = in_1265[15:0];
  assign reg_632__in[15:0] = and_632__out[15:0];
  assign and_634__in0[15:0] = in_1268[15:0];
  assign and_634__in1[15:0] = in_1269[15:0];
  assign reg_634__in[15:0] = and_634__out[15:0];
  assign and_636__in0[15:0] = in_1272[15:0];
  assign and_636__in1[15:0] = in_1273[15:0];
  assign reg_636__in[15:0] = and_636__out[15:0];
  assign and_638__in0[15:0] = in_1276[15:0];
  assign and_638__in1[15:0] = in_1277[15:0];
  assign reg_638__in[15:0] = and_638__out[15:0];
  assign and_64__in0[15:0] = in_128[15:0];
  assign and_64__in1[15:0] = in_129[15:0];
  assign reg_64__in[15:0] = and_64__out[15:0];
  assign and_640__in0[15:0] = in_1280[15:0];
  assign and_640__in1[15:0] = in_1281[15:0];
  assign reg_640__in[15:0] = and_640__out[15:0];
  assign and_642__in0[15:0] = in_1284[15:0];
  assign and_642__in1[15:0] = in_1285[15:0];
  assign reg_642__in[15:0] = and_642__out[15:0];
  assign and_644__in0[15:0] = in_1288[15:0];
  assign and_644__in1[15:0] = in_1289[15:0];
  assign reg_644__in[15:0] = and_644__out[15:0];
  assign and_646__in0[15:0] = in_1292[15:0];
  assign and_646__in1[15:0] = in_1293[15:0];
  assign reg_646__in[15:0] = and_646__out[15:0];
  assign and_648__in0[15:0] = in_1296[15:0];
  assign and_648__in1[15:0] = in_1297[15:0];
  assign reg_648__in[15:0] = and_648__out[15:0];
  assign and_650__in0[15:0] = in_1300[15:0];
  assign and_650__in1[15:0] = in_1301[15:0];
  assign reg_650__in[15:0] = and_650__out[15:0];
  assign and_652__in0[15:0] = in_1304[15:0];
  assign and_652__in1[15:0] = in_1305[15:0];
  assign reg_652__in[15:0] = and_652__out[15:0];
  assign and_654__in0[15:0] = in_1308[15:0];
  assign and_654__in1[15:0] = in_1309[15:0];
  assign reg_654__in[15:0] = and_654__out[15:0];
  assign and_656__in0[15:0] = in_1312[15:0];
  assign and_656__in1[15:0] = in_1313[15:0];
  assign reg_656__in[15:0] = and_656__out[15:0];
  assign and_658__in0[15:0] = in_1316[15:0];
  assign and_658__in1[15:0] = in_1317[15:0];
  assign reg_658__in[15:0] = and_658__out[15:0];
  assign and_66__in0[15:0] = in_132[15:0];
  assign and_66__in1[15:0] = in_133[15:0];
  assign reg_66__in[15:0] = and_66__out[15:0];
  assign and_660__in0[15:0] = in_1320[15:0];
  assign and_660__in1[15:0] = in_1321[15:0];
  assign reg_660__in[15:0] = and_660__out[15:0];
  assign and_662__in0[15:0] = in_1324[15:0];
  assign and_662__in1[15:0] = in_1325[15:0];
  assign reg_662__in[15:0] = and_662__out[15:0];
  assign and_664__in0[15:0] = in_1328[15:0];
  assign and_664__in1[15:0] = in_1329[15:0];
  assign reg_664__in[15:0] = and_664__out[15:0];
  assign and_666__in0[15:0] = in_1332[15:0];
  assign and_666__in1[15:0] = in_1333[15:0];
  assign reg_666__in[15:0] = and_666__out[15:0];
  assign and_668__in0[15:0] = in_1336[15:0];
  assign and_668__in1[15:0] = in_1337[15:0];
  assign reg_668__in[15:0] = and_668__out[15:0];
  assign and_670__in0[15:0] = in_1340[15:0];
  assign and_670__in1[15:0] = in_1341[15:0];
  assign reg_670__in[15:0] = and_670__out[15:0];
  assign and_672__in0[15:0] = in_1344[15:0];
  assign and_672__in1[15:0] = in_1345[15:0];
  assign reg_672__in[15:0] = and_672__out[15:0];
  assign and_674__in0[15:0] = in_1348[15:0];
  assign and_674__in1[15:0] = in_1349[15:0];
  assign reg_674__in[15:0] = and_674__out[15:0];
  assign and_676__in0[15:0] = in_1352[15:0];
  assign and_676__in1[15:0] = in_1353[15:0];
  assign reg_676__in[15:0] = and_676__out[15:0];
  assign and_678__in0[15:0] = in_1356[15:0];
  assign and_678__in1[15:0] = in_1357[15:0];
  assign reg_678__in[15:0] = and_678__out[15:0];
  assign and_68__in0[15:0] = in_136[15:0];
  assign and_68__in1[15:0] = in_137[15:0];
  assign reg_68__in[15:0] = and_68__out[15:0];
  assign and_680__in0[15:0] = in_1360[15:0];
  assign and_680__in1[15:0] = in_1361[15:0];
  assign reg_680__in[15:0] = and_680__out[15:0];
  assign and_682__in0[15:0] = in_1364[15:0];
  assign and_682__in1[15:0] = in_1365[15:0];
  assign reg_682__in[15:0] = and_682__out[15:0];
  assign and_684__in0[15:0] = in_1368[15:0];
  assign and_684__in1[15:0] = in_1369[15:0];
  assign reg_684__in[15:0] = and_684__out[15:0];
  assign and_686__in0[15:0] = in_1372[15:0];
  assign and_686__in1[15:0] = in_1373[15:0];
  assign reg_686__in[15:0] = and_686__out[15:0];
  assign and_688__in0[15:0] = in_1376[15:0];
  assign and_688__in1[15:0] = in_1377[15:0];
  assign reg_688__in[15:0] = and_688__out[15:0];
  assign and_690__in0[15:0] = in_1380[15:0];
  assign and_690__in1[15:0] = in_1381[15:0];
  assign reg_690__in[15:0] = and_690__out[15:0];
  assign and_692__in0[15:0] = in_1384[15:0];
  assign and_692__in1[15:0] = in_1385[15:0];
  assign reg_692__in[15:0] = and_692__out[15:0];
  assign and_694__in0[15:0] = in_1388[15:0];
  assign and_694__in1[15:0] = in_1389[15:0];
  assign reg_694__in[15:0] = and_694__out[15:0];
  assign and_696__in0[15:0] = in_1392[15:0];
  assign and_696__in1[15:0] = in_1393[15:0];
  assign reg_696__in[15:0] = and_696__out[15:0];
  assign and_698__in0[15:0] = in_1396[15:0];
  assign and_698__in1[15:0] = in_1397[15:0];
  assign reg_698__in[15:0] = and_698__out[15:0];
  assign and_70__in0[15:0] = in_140[15:0];
  assign and_70__in1[15:0] = in_141[15:0];
  assign reg_70__in[15:0] = and_70__out[15:0];
  assign and_700__in0[15:0] = in_1400[15:0];
  assign and_700__in1[15:0] = in_1401[15:0];
  assign reg_700__in[15:0] = and_700__out[15:0];
  assign and_702__in0[15:0] = in_1404[15:0];
  assign and_702__in1[15:0] = in_1405[15:0];
  assign reg_702__in[15:0] = and_702__out[15:0];
  assign and_704__in0[15:0] = in_1408[15:0];
  assign and_704__in1[15:0] = in_1409[15:0];
  assign reg_704__in[15:0] = and_704__out[15:0];
  assign and_706__in0[15:0] = in_1412[15:0];
  assign and_706__in1[15:0] = in_1413[15:0];
  assign reg_706__in[15:0] = and_706__out[15:0];
  assign and_708__in0[15:0] = in_1416[15:0];
  assign and_708__in1[15:0] = in_1417[15:0];
  assign reg_708__in[15:0] = and_708__out[15:0];
  assign and_710__in0[15:0] = in_1420[15:0];
  assign and_710__in1[15:0] = in_1421[15:0];
  assign reg_710__in[15:0] = and_710__out[15:0];
  assign and_712__in0[15:0] = in_1424[15:0];
  assign and_712__in1[15:0] = in_1425[15:0];
  assign reg_712__in[15:0] = and_712__out[15:0];
  assign and_714__in0[15:0] = in_1428[15:0];
  assign and_714__in1[15:0] = in_1429[15:0];
  assign reg_714__in[15:0] = and_714__out[15:0];
  assign and_716__in0[15:0] = in_1432[15:0];
  assign and_716__in1[15:0] = in_1433[15:0];
  assign reg_716__in[15:0] = and_716__out[15:0];
  assign and_718__in0[15:0] = in_1436[15:0];
  assign and_718__in1[15:0] = in_1437[15:0];
  assign reg_718__in[15:0] = and_718__out[15:0];
  assign and_72__in0[15:0] = in_144[15:0];
  assign and_72__in1[15:0] = in_145[15:0];
  assign reg_72__in[15:0] = and_72__out[15:0];
  assign and_720__in0[15:0] = in_1440[15:0];
  assign and_720__in1[15:0] = in_1441[15:0];
  assign reg_720__in[15:0] = and_720__out[15:0];
  assign and_722__in0[15:0] = in_1444[15:0];
  assign and_722__in1[15:0] = in_1445[15:0];
  assign reg_722__in[15:0] = and_722__out[15:0];
  assign and_724__in0[15:0] = in_1448[15:0];
  assign and_724__in1[15:0] = in_1449[15:0];
  assign reg_724__in[15:0] = and_724__out[15:0];
  assign and_726__in0[15:0] = in_1452[15:0];
  assign and_726__in1[15:0] = in_1453[15:0];
  assign reg_726__in[15:0] = and_726__out[15:0];
  assign and_728__in0[15:0] = in_1456[15:0];
  assign and_728__in1[15:0] = in_1457[15:0];
  assign reg_728__in[15:0] = and_728__out[15:0];
  assign and_730__in0[15:0] = in_1460[15:0];
  assign and_730__in1[15:0] = in_1461[15:0];
  assign reg_730__in[15:0] = and_730__out[15:0];
  assign and_732__in0[15:0] = in_1464[15:0];
  assign and_732__in1[15:0] = in_1465[15:0];
  assign reg_732__in[15:0] = and_732__out[15:0];
  assign and_734__in0[15:0] = in_1468[15:0];
  assign and_734__in1[15:0] = in_1469[15:0];
  assign reg_734__in[15:0] = and_734__out[15:0];
  assign and_736__in0[15:0] = in_1472[15:0];
  assign and_736__in1[15:0] = in_1473[15:0];
  assign reg_736__in[15:0] = and_736__out[15:0];
  assign and_738__in0[15:0] = in_1476[15:0];
  assign and_738__in1[15:0] = in_1477[15:0];
  assign reg_738__in[15:0] = and_738__out[15:0];
  assign and_74__in0[15:0] = in_148[15:0];
  assign and_74__in1[15:0] = in_149[15:0];
  assign reg_74__in[15:0] = and_74__out[15:0];
  assign and_740__in0[15:0] = in_1480[15:0];
  assign and_740__in1[15:0] = in_1481[15:0];
  assign reg_740__in[15:0] = and_740__out[15:0];
  assign and_742__in0[15:0] = in_1484[15:0];
  assign and_742__in1[15:0] = in_1485[15:0];
  assign reg_742__in[15:0] = and_742__out[15:0];
  assign and_744__in0[15:0] = in_1488[15:0];
  assign and_744__in1[15:0] = in_1489[15:0];
  assign reg_744__in[15:0] = and_744__out[15:0];
  assign and_746__in0[15:0] = in_1492[15:0];
  assign and_746__in1[15:0] = in_1493[15:0];
  assign reg_746__in[15:0] = and_746__out[15:0];
  assign and_748__in0[15:0] = in_1496[15:0];
  assign and_748__in1[15:0] = in_1497[15:0];
  assign reg_748__in[15:0] = and_748__out[15:0];
  assign and_750__in0[15:0] = in_1500[15:0];
  assign and_750__in1[15:0] = in_1501[15:0];
  assign reg_750__in[15:0] = and_750__out[15:0];
  assign and_752__in0[15:0] = in_1504[15:0];
  assign and_752__in1[15:0] = in_1505[15:0];
  assign reg_752__in[15:0] = and_752__out[15:0];
  assign and_754__in0[15:0] = in_1508[15:0];
  assign and_754__in1[15:0] = in_1509[15:0];
  assign reg_754__in[15:0] = and_754__out[15:0];
  assign and_756__in0[15:0] = in_1512[15:0];
  assign and_756__in1[15:0] = in_1513[15:0];
  assign reg_756__in[15:0] = and_756__out[15:0];
  assign and_758__in0[15:0] = in_1516[15:0];
  assign and_758__in1[15:0] = in_1517[15:0];
  assign reg_758__in[15:0] = and_758__out[15:0];
  assign and_76__in0[15:0] = in_152[15:0];
  assign and_76__in1[15:0] = in_153[15:0];
  assign reg_76__in[15:0] = and_76__out[15:0];
  assign and_760__in0[15:0] = in_1520[15:0];
  assign and_760__in1[15:0] = in_1521[15:0];
  assign reg_760__in[15:0] = and_760__out[15:0];
  assign and_762__in0[15:0] = in_1524[15:0];
  assign and_762__in1[15:0] = in_1525[15:0];
  assign reg_762__in[15:0] = and_762__out[15:0];
  assign and_764__in0[15:0] = in_1528[15:0];
  assign and_764__in1[15:0] = in_1529[15:0];
  assign reg_764__in[15:0] = and_764__out[15:0];
  assign and_766__in0[15:0] = in_1532[15:0];
  assign and_766__in1[15:0] = in_1533[15:0];
  assign reg_766__in[15:0] = and_766__out[15:0];
  assign and_768__in0[15:0] = in_1536[15:0];
  assign and_768__in1[15:0] = in_1537[15:0];
  assign reg_768__in[15:0] = and_768__out[15:0];
  assign and_770__in0[15:0] = in_1540[15:0];
  assign and_770__in1[15:0] = in_1541[15:0];
  assign reg_770__in[15:0] = and_770__out[15:0];
  assign and_772__in0[15:0] = in_1544[15:0];
  assign and_772__in1[15:0] = in_1545[15:0];
  assign reg_772__in[15:0] = and_772__out[15:0];
  assign and_774__in0[15:0] = in_1548[15:0];
  assign and_774__in1[15:0] = in_1549[15:0];
  assign reg_774__in[15:0] = and_774__out[15:0];
  assign and_776__in0[15:0] = in_1552[15:0];
  assign and_776__in1[15:0] = in_1553[15:0];
  assign reg_776__in[15:0] = and_776__out[15:0];
  assign and_778__in0[15:0] = in_1556[15:0];
  assign and_778__in1[15:0] = in_1557[15:0];
  assign reg_778__in[15:0] = and_778__out[15:0];
  assign and_78__in0[15:0] = in_156[15:0];
  assign and_78__in1[15:0] = in_157[15:0];
  assign reg_78__in[15:0] = and_78__out[15:0];
  assign and_780__in0[15:0] = in_1560[15:0];
  assign and_780__in1[15:0] = in_1561[15:0];
  assign reg_780__in[15:0] = and_780__out[15:0];
  assign and_782__in0[15:0] = in_1564[15:0];
  assign and_782__in1[15:0] = in_1565[15:0];
  assign reg_782__in[15:0] = and_782__out[15:0];
  assign and_784__in0[15:0] = in_1568[15:0];
  assign and_784__in1[15:0] = in_1569[15:0];
  assign reg_784__in[15:0] = and_784__out[15:0];
  assign and_786__in0[15:0] = in_1572[15:0];
  assign and_786__in1[15:0] = in_1573[15:0];
  assign reg_786__in[15:0] = and_786__out[15:0];
  assign and_788__in0[15:0] = in_1576[15:0];
  assign and_788__in1[15:0] = in_1577[15:0];
  assign reg_788__in[15:0] = and_788__out[15:0];
  assign and_790__in0[15:0] = in_1580[15:0];
  assign and_790__in1[15:0] = in_1581[15:0];
  assign reg_790__in[15:0] = and_790__out[15:0];
  assign and_792__in0[15:0] = in_1584[15:0];
  assign and_792__in1[15:0] = in_1585[15:0];
  assign reg_792__in[15:0] = and_792__out[15:0];
  assign and_794__in0[15:0] = in_1588[15:0];
  assign and_794__in1[15:0] = in_1589[15:0];
  assign reg_794__in[15:0] = and_794__out[15:0];
  assign and_796__in0[15:0] = in_1592[15:0];
  assign and_796__in1[15:0] = in_1593[15:0];
  assign reg_796__in[15:0] = and_796__out[15:0];
  assign and_798__in0[15:0] = in_1596[15:0];
  assign and_798__in1[15:0] = in_1597[15:0];
  assign reg_798__in[15:0] = and_798__out[15:0];
  assign and_8__in0[15:0] = in_16[15:0];
  assign and_8__in1[15:0] = in_17[15:0];
  assign reg_8__in[15:0] = and_8__out[15:0];
  assign and_80__in0[15:0] = in_160[15:0];
  assign and_80__in1[15:0] = in_161[15:0];
  assign reg_80__in[15:0] = and_80__out[15:0];
  assign and_800__in0[15:0] = in_1600[15:0];
  assign and_800__in1[15:0] = in_1601[15:0];
  assign reg_800__in[15:0] = and_800__out[15:0];
  assign and_802__in0[15:0] = in_1604[15:0];
  assign and_802__in1[15:0] = in_1605[15:0];
  assign reg_802__in[15:0] = and_802__out[15:0];
  assign and_804__in0[15:0] = in_1608[15:0];
  assign and_804__in1[15:0] = in_1609[15:0];
  assign reg_804__in[15:0] = and_804__out[15:0];
  assign and_806__in0[15:0] = in_1612[15:0];
  assign and_806__in1[15:0] = in_1613[15:0];
  assign reg_806__in[15:0] = and_806__out[15:0];
  assign and_808__in0[15:0] = in_1616[15:0];
  assign and_808__in1[15:0] = in_1617[15:0];
  assign reg_808__in[15:0] = and_808__out[15:0];
  assign and_810__in0[15:0] = in_1620[15:0];
  assign and_810__in1[15:0] = in_1621[15:0];
  assign reg_810__in[15:0] = and_810__out[15:0];
  assign and_812__in0[15:0] = in_1624[15:0];
  assign and_812__in1[15:0] = in_1625[15:0];
  assign reg_812__in[15:0] = and_812__out[15:0];
  assign and_814__in0[15:0] = in_1628[15:0];
  assign and_814__in1[15:0] = in_1629[15:0];
  assign reg_814__in[15:0] = and_814__out[15:0];
  assign and_816__in0[15:0] = in_1632[15:0];
  assign and_816__in1[15:0] = in_1633[15:0];
  assign reg_816__in[15:0] = and_816__out[15:0];
  assign and_818__in0[15:0] = in_1636[15:0];
  assign and_818__in1[15:0] = in_1637[15:0];
  assign reg_818__in[15:0] = and_818__out[15:0];
  assign and_82__in0[15:0] = in_164[15:0];
  assign and_82__in1[15:0] = in_165[15:0];
  assign reg_82__in[15:0] = and_82__out[15:0];
  assign and_820__in0[15:0] = in_1640[15:0];
  assign and_820__in1[15:0] = in_1641[15:0];
  assign reg_820__in[15:0] = and_820__out[15:0];
  assign and_822__in0[15:0] = in_1644[15:0];
  assign and_822__in1[15:0] = in_1645[15:0];
  assign reg_822__in[15:0] = and_822__out[15:0];
  assign and_824__in0[15:0] = in_1648[15:0];
  assign and_824__in1[15:0] = in_1649[15:0];
  assign reg_824__in[15:0] = and_824__out[15:0];
  assign and_826__in0[15:0] = in_1652[15:0];
  assign and_826__in1[15:0] = in_1653[15:0];
  assign reg_826__in[15:0] = and_826__out[15:0];
  assign and_828__in0[15:0] = in_1656[15:0];
  assign and_828__in1[15:0] = in_1657[15:0];
  assign reg_828__in[15:0] = and_828__out[15:0];
  assign and_830__in0[15:0] = in_1660[15:0];
  assign and_830__in1[15:0] = in_1661[15:0];
  assign reg_830__in[15:0] = and_830__out[15:0];
  assign and_832__in0[15:0] = in_1664[15:0];
  assign and_832__in1[15:0] = in_1665[15:0];
  assign reg_832__in[15:0] = and_832__out[15:0];
  assign and_834__in0[15:0] = in_1668[15:0];
  assign and_834__in1[15:0] = in_1669[15:0];
  assign reg_834__in[15:0] = and_834__out[15:0];
  assign and_836__in0[15:0] = in_1672[15:0];
  assign and_836__in1[15:0] = in_1673[15:0];
  assign reg_836__in[15:0] = and_836__out[15:0];
  assign and_838__in0[15:0] = in_1676[15:0];
  assign and_838__in1[15:0] = in_1677[15:0];
  assign reg_838__in[15:0] = and_838__out[15:0];
  assign and_84__in0[15:0] = in_168[15:0];
  assign and_84__in1[15:0] = in_169[15:0];
  assign reg_84__in[15:0] = and_84__out[15:0];
  assign and_840__in0[15:0] = in_1680[15:0];
  assign and_840__in1[15:0] = in_1681[15:0];
  assign reg_840__in[15:0] = and_840__out[15:0];
  assign and_842__in0[15:0] = in_1684[15:0];
  assign and_842__in1[15:0] = in_1685[15:0];
  assign reg_842__in[15:0] = and_842__out[15:0];
  assign and_844__in0[15:0] = in_1688[15:0];
  assign and_844__in1[15:0] = in_1689[15:0];
  assign reg_844__in[15:0] = and_844__out[15:0];
  assign and_846__in0[15:0] = in_1692[15:0];
  assign and_846__in1[15:0] = in_1693[15:0];
  assign reg_846__in[15:0] = and_846__out[15:0];
  assign and_848__in0[15:0] = in_1696[15:0];
  assign and_848__in1[15:0] = in_1697[15:0];
  assign reg_848__in[15:0] = and_848__out[15:0];
  assign and_850__in0[15:0] = in_1700[15:0];
  assign and_850__in1[15:0] = in_1701[15:0];
  assign reg_850__in[15:0] = and_850__out[15:0];
  assign and_852__in0[15:0] = in_1704[15:0];
  assign and_852__in1[15:0] = in_1705[15:0];
  assign reg_852__in[15:0] = and_852__out[15:0];
  assign and_854__in0[15:0] = in_1708[15:0];
  assign and_854__in1[15:0] = in_1709[15:0];
  assign reg_854__in[15:0] = and_854__out[15:0];
  assign and_856__in0[15:0] = in_1712[15:0];
  assign and_856__in1[15:0] = in_1713[15:0];
  assign reg_856__in[15:0] = and_856__out[15:0];
  assign and_858__in0[15:0] = in_1716[15:0];
  assign and_858__in1[15:0] = in_1717[15:0];
  assign reg_858__in[15:0] = and_858__out[15:0];
  assign and_86__in0[15:0] = in_172[15:0];
  assign and_86__in1[15:0] = in_173[15:0];
  assign reg_86__in[15:0] = and_86__out[15:0];
  assign and_860__in0[15:0] = in_1720[15:0];
  assign and_860__in1[15:0] = in_1721[15:0];
  assign reg_860__in[15:0] = and_860__out[15:0];
  assign and_862__in0[15:0] = in_1724[15:0];
  assign and_862__in1[15:0] = in_1725[15:0];
  assign reg_862__in[15:0] = and_862__out[15:0];
  assign and_864__in0[15:0] = in_1728[15:0];
  assign and_864__in1[15:0] = in_1729[15:0];
  assign reg_864__in[15:0] = and_864__out[15:0];
  assign and_866__in0[15:0] = in_1732[15:0];
  assign and_866__in1[15:0] = in_1733[15:0];
  assign reg_866__in[15:0] = and_866__out[15:0];
  assign and_868__in0[15:0] = in_1736[15:0];
  assign and_868__in1[15:0] = in_1737[15:0];
  assign reg_868__in[15:0] = and_868__out[15:0];
  assign and_870__in0[15:0] = in_1740[15:0];
  assign and_870__in1[15:0] = in_1741[15:0];
  assign reg_870__in[15:0] = and_870__out[15:0];
  assign and_872__in0[15:0] = in_1744[15:0];
  assign and_872__in1[15:0] = in_1745[15:0];
  assign reg_872__in[15:0] = and_872__out[15:0];
  assign and_874__in0[15:0] = in_1748[15:0];
  assign and_874__in1[15:0] = in_1749[15:0];
  assign reg_874__in[15:0] = and_874__out[15:0];
  assign and_876__in0[15:0] = in_1752[15:0];
  assign and_876__in1[15:0] = in_1753[15:0];
  assign reg_876__in[15:0] = and_876__out[15:0];
  assign and_878__in0[15:0] = in_1756[15:0];
  assign and_878__in1[15:0] = in_1757[15:0];
  assign reg_878__in[15:0] = and_878__out[15:0];
  assign and_88__in0[15:0] = in_176[15:0];
  assign and_88__in1[15:0] = in_177[15:0];
  assign reg_88__in[15:0] = and_88__out[15:0];
  assign and_880__in0[15:0] = in_1760[15:0];
  assign and_880__in1[15:0] = in_1761[15:0];
  assign reg_880__in[15:0] = and_880__out[15:0];
  assign and_882__in0[15:0] = in_1764[15:0];
  assign and_882__in1[15:0] = in_1765[15:0];
  assign reg_882__in[15:0] = and_882__out[15:0];
  assign and_884__in0[15:0] = in_1768[15:0];
  assign and_884__in1[15:0] = in_1769[15:0];
  assign reg_884__in[15:0] = and_884__out[15:0];
  assign and_886__in0[15:0] = in_1772[15:0];
  assign and_886__in1[15:0] = in_1773[15:0];
  assign reg_886__in[15:0] = and_886__out[15:0];
  assign and_888__in0[15:0] = in_1776[15:0];
  assign and_888__in1[15:0] = in_1777[15:0];
  assign reg_888__in[15:0] = and_888__out[15:0];
  assign and_890__in0[15:0] = in_1780[15:0];
  assign and_890__in1[15:0] = in_1781[15:0];
  assign reg_890__in[15:0] = and_890__out[15:0];
  assign and_892__in0[15:0] = in_1784[15:0];
  assign and_892__in1[15:0] = in_1785[15:0];
  assign reg_892__in[15:0] = and_892__out[15:0];
  assign and_894__in0[15:0] = in_1788[15:0];
  assign and_894__in1[15:0] = in_1789[15:0];
  assign reg_894__in[15:0] = and_894__out[15:0];
  assign and_896__in0[15:0] = in_1792[15:0];
  assign and_896__in1[15:0] = in_1793[15:0];
  assign reg_896__in[15:0] = and_896__out[15:0];
  assign and_898__in0[15:0] = in_1796[15:0];
  assign and_898__in1[15:0] = in_1797[15:0];
  assign reg_898__in[15:0] = and_898__out[15:0];
  assign and_90__in0[15:0] = in_180[15:0];
  assign and_90__in1[15:0] = in_181[15:0];
  assign reg_90__in[15:0] = and_90__out[15:0];
  assign and_900__in0[15:0] = in_1800[15:0];
  assign and_900__in1[15:0] = in_1801[15:0];
  assign reg_900__in[15:0] = and_900__out[15:0];
  assign and_902__in0[15:0] = in_1804[15:0];
  assign and_902__in1[15:0] = in_1805[15:0];
  assign reg_902__in[15:0] = and_902__out[15:0];
  assign and_904__in0[15:0] = in_1808[15:0];
  assign and_904__in1[15:0] = in_1809[15:0];
  assign reg_904__in[15:0] = and_904__out[15:0];
  assign and_906__in0[15:0] = in_1812[15:0];
  assign and_906__in1[15:0] = in_1813[15:0];
  assign reg_906__in[15:0] = and_906__out[15:0];
  assign and_908__in0[15:0] = in_1816[15:0];
  assign and_908__in1[15:0] = in_1817[15:0];
  assign reg_908__in[15:0] = and_908__out[15:0];
  assign and_910__in0[15:0] = in_1820[15:0];
  assign and_910__in1[15:0] = in_1821[15:0];
  assign reg_910__in[15:0] = and_910__out[15:0];
  assign and_912__in0[15:0] = in_1824[15:0];
  assign and_912__in1[15:0] = in_1825[15:0];
  assign reg_912__in[15:0] = and_912__out[15:0];
  assign and_914__in0[15:0] = in_1828[15:0];
  assign and_914__in1[15:0] = in_1829[15:0];
  assign reg_914__in[15:0] = and_914__out[15:0];
  assign and_916__in0[15:0] = in_1832[15:0];
  assign and_916__in1[15:0] = in_1833[15:0];
  assign reg_916__in[15:0] = and_916__out[15:0];
  assign and_918__in0[15:0] = in_1836[15:0];
  assign and_918__in1[15:0] = in_1837[15:0];
  assign reg_918__in[15:0] = and_918__out[15:0];
  assign and_92__in0[15:0] = in_184[15:0];
  assign and_92__in1[15:0] = in_185[15:0];
  assign reg_92__in[15:0] = and_92__out[15:0];
  assign and_920__in0[15:0] = in_1840[15:0];
  assign and_920__in1[15:0] = in_1841[15:0];
  assign reg_920__in[15:0] = and_920__out[15:0];
  assign and_922__in0[15:0] = in_1844[15:0];
  assign and_922__in1[15:0] = in_1845[15:0];
  assign reg_922__in[15:0] = and_922__out[15:0];
  assign and_924__in0[15:0] = in_1848[15:0];
  assign and_924__in1[15:0] = in_1849[15:0];
  assign reg_924__in[15:0] = and_924__out[15:0];
  assign and_926__in0[15:0] = in_1852[15:0];
  assign and_926__in1[15:0] = in_1853[15:0];
  assign reg_926__in[15:0] = and_926__out[15:0];
  assign and_928__in0[15:0] = in_1856[15:0];
  assign and_928__in1[15:0] = in_1857[15:0];
  assign reg_928__in[15:0] = and_928__out[15:0];
  assign and_930__in0[15:0] = in_1860[15:0];
  assign and_930__in1[15:0] = in_1861[15:0];
  assign reg_930__in[15:0] = and_930__out[15:0];
  assign and_932__in0[15:0] = in_1864[15:0];
  assign and_932__in1[15:0] = in_1865[15:0];
  assign reg_932__in[15:0] = and_932__out[15:0];
  assign and_934__in0[15:0] = in_1868[15:0];
  assign and_934__in1[15:0] = in_1869[15:0];
  assign reg_934__in[15:0] = and_934__out[15:0];
  assign and_936__in0[15:0] = in_1872[15:0];
  assign and_936__in1[15:0] = in_1873[15:0];
  assign reg_936__in[15:0] = and_936__out[15:0];
  assign and_938__in0[15:0] = in_1876[15:0];
  assign and_938__in1[15:0] = in_1877[15:0];
  assign reg_938__in[15:0] = and_938__out[15:0];
  assign and_94__in0[15:0] = in_188[15:0];
  assign and_94__in1[15:0] = in_189[15:0];
  assign reg_94__in[15:0] = and_94__out[15:0];
  assign and_940__in0[15:0] = in_1880[15:0];
  assign and_940__in1[15:0] = in_1881[15:0];
  assign reg_940__in[15:0] = and_940__out[15:0];
  assign and_942__in0[15:0] = in_1884[15:0];
  assign and_942__in1[15:0] = in_1885[15:0];
  assign reg_942__in[15:0] = and_942__out[15:0];
  assign and_944__in0[15:0] = in_1888[15:0];
  assign and_944__in1[15:0] = in_1889[15:0];
  assign reg_944__in[15:0] = and_944__out[15:0];
  assign and_946__in0[15:0] = in_1892[15:0];
  assign and_946__in1[15:0] = in_1893[15:0];
  assign reg_946__in[15:0] = and_946__out[15:0];
  assign and_948__in0[15:0] = in_1896[15:0];
  assign and_948__in1[15:0] = in_1897[15:0];
  assign reg_948__in[15:0] = and_948__out[15:0];
  assign and_950__in0[15:0] = in_1900[15:0];
  assign and_950__in1[15:0] = in_1901[15:0];
  assign reg_950__in[15:0] = and_950__out[15:0];
  assign and_952__in0[15:0] = in_1904[15:0];
  assign and_952__in1[15:0] = in_1905[15:0];
  assign reg_952__in[15:0] = and_952__out[15:0];
  assign and_954__in0[15:0] = in_1908[15:0];
  assign and_954__in1[15:0] = in_1909[15:0];
  assign reg_954__in[15:0] = and_954__out[15:0];
  assign and_956__in0[15:0] = in_1912[15:0];
  assign and_956__in1[15:0] = in_1913[15:0];
  assign reg_956__in[15:0] = and_956__out[15:0];
  assign and_958__in0[15:0] = in_1916[15:0];
  assign and_958__in1[15:0] = in_1917[15:0];
  assign reg_958__in[15:0] = and_958__out[15:0];
  assign and_96__in0[15:0] = in_192[15:0];
  assign and_96__in1[15:0] = in_193[15:0];
  assign reg_96__in[15:0] = and_96__out[15:0];
  assign and_960__in0[15:0] = in_1920[15:0];
  assign and_960__in1[15:0] = in_1921[15:0];
  assign reg_960__in[15:0] = and_960__out[15:0];
  assign and_962__in0[15:0] = in_1924[15:0];
  assign and_962__in1[15:0] = in_1925[15:0];
  assign reg_962__in[15:0] = and_962__out[15:0];
  assign and_964__in0[15:0] = in_1928[15:0];
  assign and_964__in1[15:0] = in_1929[15:0];
  assign reg_964__in[15:0] = and_964__out[15:0];
  assign and_966__in0[15:0] = in_1932[15:0];
  assign and_966__in1[15:0] = in_1933[15:0];
  assign reg_966__in[15:0] = and_966__out[15:0];
  assign and_968__in0[15:0] = in_1936[15:0];
  assign and_968__in1[15:0] = in_1937[15:0];
  assign reg_968__in[15:0] = and_968__out[15:0];
  assign and_970__in0[15:0] = in_1940[15:0];
  assign and_970__in1[15:0] = in_1941[15:0];
  assign reg_970__in[15:0] = and_970__out[15:0];
  assign and_972__in0[15:0] = in_1944[15:0];
  assign and_972__in1[15:0] = in_1945[15:0];
  assign reg_972__in[15:0] = and_972__out[15:0];
  assign and_974__in0[15:0] = in_1948[15:0];
  assign and_974__in1[15:0] = in_1949[15:0];
  assign reg_974__in[15:0] = and_974__out[15:0];
  assign and_976__in0[15:0] = in_1952[15:0];
  assign and_976__in1[15:0] = in_1953[15:0];
  assign reg_976__in[15:0] = and_976__out[15:0];
  assign and_978__in0[15:0] = in_1956[15:0];
  assign and_978__in1[15:0] = in_1957[15:0];
  assign reg_978__in[15:0] = and_978__out[15:0];
  assign and_98__in0[15:0] = in_196[15:0];
  assign and_98__in1[15:0] = in_197[15:0];
  assign reg_98__in[15:0] = and_98__out[15:0];
  assign and_980__in0[15:0] = in_1960[15:0];
  assign and_980__in1[15:0] = in_1961[15:0];
  assign reg_980__in[15:0] = and_980__out[15:0];
  assign and_982__in0[15:0] = in_1964[15:0];
  assign and_982__in1[15:0] = in_1965[15:0];
  assign reg_982__in[15:0] = and_982__out[15:0];
  assign and_984__in0[15:0] = in_1968[15:0];
  assign and_984__in1[15:0] = in_1969[15:0];
  assign reg_984__in[15:0] = and_984__out[15:0];
  assign and_986__in0[15:0] = in_1972[15:0];
  assign and_986__in1[15:0] = in_1973[15:0];
  assign reg_986__in[15:0] = and_986__out[15:0];
  assign and_988__in0[15:0] = in_1976[15:0];
  assign and_988__in1[15:0] = in_1977[15:0];
  assign reg_988__in[15:0] = and_988__out[15:0];
  assign and_990__in0[15:0] = in_1980[15:0];
  assign and_990__in1[15:0] = in_1981[15:0];
  assign reg_990__in[15:0] = and_990__out[15:0];
  assign and_992__in0[15:0] = in_1984[15:0];
  assign and_992__in1[15:0] = in_1985[15:0];
  assign reg_992__in[15:0] = and_992__out[15:0];
  assign and_994__in0[15:0] = in_1988[15:0];
  assign and_994__in1[15:0] = in_1989[15:0];
  assign reg_994__in[15:0] = and_994__out[15:0];
  assign and_996__in0[15:0] = in_1992[15:0];
  assign and_996__in1[15:0] = in_1993[15:0];
  assign reg_996__in[15:0] = and_996__out[15:0];
  assign and_998__in0[15:0] = in_1996[15:0];
  assign and_998__in1[15:0] = in_1997[15:0];
  assign reg_998__in[15:0] = and_998__out[15:0];
  assign or_1__in0[15:0] = in_2[15:0];
  assign or_1__in1[15:0] = in_3[15:0];
  assign reg_1__in[15:0] = or_1__out[15:0];
  assign or_101__in0[15:0] = in_202[15:0];
  assign or_101__in1[15:0] = in_203[15:0];
  assign reg_101__in[15:0] = or_101__out[15:0];
  assign or_103__in0[15:0] = in_206[15:0];
  assign or_103__in1[15:0] = in_207[15:0];
  assign reg_103__in[15:0] = or_103__out[15:0];
  assign or_105__in0[15:0] = in_210[15:0];
  assign or_105__in1[15:0] = in_211[15:0];
  assign reg_105__in[15:0] = or_105__out[15:0];
  assign or_107__in0[15:0] = in_214[15:0];
  assign or_107__in1[15:0] = in_215[15:0];
  assign reg_107__in[15:0] = or_107__out[15:0];
  assign or_109__in0[15:0] = in_218[15:0];
  assign or_109__in1[15:0] = in_219[15:0];
  assign reg_109__in[15:0] = or_109__out[15:0];
  assign or_11__in0[15:0] = in_22[15:0];
  assign or_11__in1[15:0] = in_23[15:0];
  assign reg_11__in[15:0] = or_11__out[15:0];
  assign or_111__in0[15:0] = in_222[15:0];
  assign or_111__in1[15:0] = in_223[15:0];
  assign reg_111__in[15:0] = or_111__out[15:0];
  assign or_113__in0[15:0] = in_226[15:0];
  assign or_113__in1[15:0] = in_227[15:0];
  assign reg_113__in[15:0] = or_113__out[15:0];
  assign or_115__in0[15:0] = in_230[15:0];
  assign or_115__in1[15:0] = in_231[15:0];
  assign reg_115__in[15:0] = or_115__out[15:0];
  assign or_117__in0[15:0] = in_234[15:0];
  assign or_117__in1[15:0] = in_235[15:0];
  assign reg_117__in[15:0] = or_117__out[15:0];
  assign or_119__in0[15:0] = in_238[15:0];
  assign or_119__in1[15:0] = in_239[15:0];
  assign reg_119__in[15:0] = or_119__out[15:0];
  assign or_121__in0[15:0] = in_242[15:0];
  assign or_121__in1[15:0] = in_243[15:0];
  assign reg_121__in[15:0] = or_121__out[15:0];
  assign or_123__in0[15:0] = in_246[15:0];
  assign or_123__in1[15:0] = in_247[15:0];
  assign reg_123__in[15:0] = or_123__out[15:0];
  assign or_125__in0[15:0] = in_250[15:0];
  assign or_125__in1[15:0] = in_251[15:0];
  assign reg_125__in[15:0] = or_125__out[15:0];
  assign or_127__in0[15:0] = in_254[15:0];
  assign or_127__in1[15:0] = in_255[15:0];
  assign reg_127__in[15:0] = or_127__out[15:0];
  assign or_129__in0[15:0] = in_258[15:0];
  assign or_129__in1[15:0] = in_259[15:0];
  assign reg_129__in[15:0] = or_129__out[15:0];
  assign or_13__in0[15:0] = in_26[15:0];
  assign or_13__in1[15:0] = in_27[15:0];
  assign reg_13__in[15:0] = or_13__out[15:0];
  assign or_131__in0[15:0] = in_262[15:0];
  assign or_131__in1[15:0] = in_263[15:0];
  assign reg_131__in[15:0] = or_131__out[15:0];
  assign or_133__in0[15:0] = in_266[15:0];
  assign or_133__in1[15:0] = in_267[15:0];
  assign reg_133__in[15:0] = or_133__out[15:0];
  assign or_135__in0[15:0] = in_270[15:0];
  assign or_135__in1[15:0] = in_271[15:0];
  assign reg_135__in[15:0] = or_135__out[15:0];
  assign or_137__in0[15:0] = in_274[15:0];
  assign or_137__in1[15:0] = in_275[15:0];
  assign reg_137__in[15:0] = or_137__out[15:0];
  assign or_139__in0[15:0] = in_278[15:0];
  assign or_139__in1[15:0] = in_279[15:0];
  assign reg_139__in[15:0] = or_139__out[15:0];
  assign or_141__in0[15:0] = in_282[15:0];
  assign or_141__in1[15:0] = in_283[15:0];
  assign reg_141__in[15:0] = or_141__out[15:0];
  assign or_143__in0[15:0] = in_286[15:0];
  assign or_143__in1[15:0] = in_287[15:0];
  assign reg_143__in[15:0] = or_143__out[15:0];
  assign or_145__in0[15:0] = in_290[15:0];
  assign or_145__in1[15:0] = in_291[15:0];
  assign reg_145__in[15:0] = or_145__out[15:0];
  assign or_147__in0[15:0] = in_294[15:0];
  assign or_147__in1[15:0] = in_295[15:0];
  assign reg_147__in[15:0] = or_147__out[15:0];
  assign or_149__in0[15:0] = in_298[15:0];
  assign or_149__in1[15:0] = in_299[15:0];
  assign reg_149__in[15:0] = or_149__out[15:0];
  assign or_15__in0[15:0] = in_30[15:0];
  assign or_15__in1[15:0] = in_31[15:0];
  assign reg_15__in[15:0] = or_15__out[15:0];
  assign or_151__in0[15:0] = in_302[15:0];
  assign or_151__in1[15:0] = in_303[15:0];
  assign reg_151__in[15:0] = or_151__out[15:0];
  assign or_153__in0[15:0] = in_306[15:0];
  assign or_153__in1[15:0] = in_307[15:0];
  assign reg_153__in[15:0] = or_153__out[15:0];
  assign or_155__in0[15:0] = in_310[15:0];
  assign or_155__in1[15:0] = in_311[15:0];
  assign reg_155__in[15:0] = or_155__out[15:0];
  assign or_157__in0[15:0] = in_314[15:0];
  assign or_157__in1[15:0] = in_315[15:0];
  assign reg_157__in[15:0] = or_157__out[15:0];
  assign or_159__in0[15:0] = in_318[15:0];
  assign or_159__in1[15:0] = in_319[15:0];
  assign reg_159__in[15:0] = or_159__out[15:0];
  assign or_161__in0[15:0] = in_322[15:0];
  assign or_161__in1[15:0] = in_323[15:0];
  assign reg_161__in[15:0] = or_161__out[15:0];
  assign or_163__in0[15:0] = in_326[15:0];
  assign or_163__in1[15:0] = in_327[15:0];
  assign reg_163__in[15:0] = or_163__out[15:0];
  assign or_165__in0[15:0] = in_330[15:0];
  assign or_165__in1[15:0] = in_331[15:0];
  assign reg_165__in[15:0] = or_165__out[15:0];
  assign or_167__in0[15:0] = in_334[15:0];
  assign or_167__in1[15:0] = in_335[15:0];
  assign reg_167__in[15:0] = or_167__out[15:0];
  assign or_169__in0[15:0] = in_338[15:0];
  assign or_169__in1[15:0] = in_339[15:0];
  assign reg_169__in[15:0] = or_169__out[15:0];
  assign or_17__in0[15:0] = in_34[15:0];
  assign or_17__in1[15:0] = in_35[15:0];
  assign reg_17__in[15:0] = or_17__out[15:0];
  assign or_171__in0[15:0] = in_342[15:0];
  assign or_171__in1[15:0] = in_343[15:0];
  assign reg_171__in[15:0] = or_171__out[15:0];
  assign or_173__in0[15:0] = in_346[15:0];
  assign or_173__in1[15:0] = in_347[15:0];
  assign reg_173__in[15:0] = or_173__out[15:0];
  assign or_175__in0[15:0] = in_350[15:0];
  assign or_175__in1[15:0] = in_351[15:0];
  assign reg_175__in[15:0] = or_175__out[15:0];
  assign or_177__in0[15:0] = in_354[15:0];
  assign or_177__in1[15:0] = in_355[15:0];
  assign reg_177__in[15:0] = or_177__out[15:0];
  assign or_179__in0[15:0] = in_358[15:0];
  assign or_179__in1[15:0] = in_359[15:0];
  assign reg_179__in[15:0] = or_179__out[15:0];
  assign or_181__in0[15:0] = in_362[15:0];
  assign or_181__in1[15:0] = in_363[15:0];
  assign reg_181__in[15:0] = or_181__out[15:0];
  assign or_183__in0[15:0] = in_366[15:0];
  assign or_183__in1[15:0] = in_367[15:0];
  assign reg_183__in[15:0] = or_183__out[15:0];
  assign or_185__in0[15:0] = in_370[15:0];
  assign or_185__in1[15:0] = in_371[15:0];
  assign reg_185__in[15:0] = or_185__out[15:0];
  assign or_187__in0[15:0] = in_374[15:0];
  assign or_187__in1[15:0] = in_375[15:0];
  assign reg_187__in[15:0] = or_187__out[15:0];
  assign or_189__in0[15:0] = in_378[15:0];
  assign or_189__in1[15:0] = in_379[15:0];
  assign reg_189__in[15:0] = or_189__out[15:0];
  assign or_19__in0[15:0] = in_38[15:0];
  assign or_19__in1[15:0] = in_39[15:0];
  assign reg_19__in[15:0] = or_19__out[15:0];
  assign or_191__in0[15:0] = in_382[15:0];
  assign or_191__in1[15:0] = in_383[15:0];
  assign reg_191__in[15:0] = or_191__out[15:0];
  assign or_193__in0[15:0] = in_386[15:0];
  assign or_193__in1[15:0] = in_387[15:0];
  assign reg_193__in[15:0] = or_193__out[15:0];
  assign or_195__in0[15:0] = in_390[15:0];
  assign or_195__in1[15:0] = in_391[15:0];
  assign reg_195__in[15:0] = or_195__out[15:0];
  assign or_197__in0[15:0] = in_394[15:0];
  assign or_197__in1[15:0] = in_395[15:0];
  assign reg_197__in[15:0] = or_197__out[15:0];
  assign or_199__in0[15:0] = in_398[15:0];
  assign or_199__in1[15:0] = in_399[15:0];
  assign reg_199__in[15:0] = or_199__out[15:0];
  assign or_201__in0[15:0] = in_402[15:0];
  assign or_201__in1[15:0] = in_403[15:0];
  assign reg_201__in[15:0] = or_201__out[15:0];
  assign or_203__in0[15:0] = in_406[15:0];
  assign or_203__in1[15:0] = in_407[15:0];
  assign reg_203__in[15:0] = or_203__out[15:0];
  assign or_205__in0[15:0] = in_410[15:0];
  assign or_205__in1[15:0] = in_411[15:0];
  assign reg_205__in[15:0] = or_205__out[15:0];
  assign or_207__in0[15:0] = in_414[15:0];
  assign or_207__in1[15:0] = in_415[15:0];
  assign reg_207__in[15:0] = or_207__out[15:0];
  assign or_209__in0[15:0] = in_418[15:0];
  assign or_209__in1[15:0] = in_419[15:0];
  assign reg_209__in[15:0] = or_209__out[15:0];
  assign or_21__in0[15:0] = in_42[15:0];
  assign or_21__in1[15:0] = in_43[15:0];
  assign reg_21__in[15:0] = or_21__out[15:0];
  assign or_211__in0[15:0] = in_422[15:0];
  assign or_211__in1[15:0] = in_423[15:0];
  assign reg_211__in[15:0] = or_211__out[15:0];
  assign or_213__in0[15:0] = in_426[15:0];
  assign or_213__in1[15:0] = in_427[15:0];
  assign reg_213__in[15:0] = or_213__out[15:0];
  assign or_215__in0[15:0] = in_430[15:0];
  assign or_215__in1[15:0] = in_431[15:0];
  assign reg_215__in[15:0] = or_215__out[15:0];
  assign or_217__in0[15:0] = in_434[15:0];
  assign or_217__in1[15:0] = in_435[15:0];
  assign reg_217__in[15:0] = or_217__out[15:0];
  assign or_219__in0[15:0] = in_438[15:0];
  assign or_219__in1[15:0] = in_439[15:0];
  assign reg_219__in[15:0] = or_219__out[15:0];
  assign or_221__in0[15:0] = in_442[15:0];
  assign or_221__in1[15:0] = in_443[15:0];
  assign reg_221__in[15:0] = or_221__out[15:0];
  assign or_223__in0[15:0] = in_446[15:0];
  assign or_223__in1[15:0] = in_447[15:0];
  assign reg_223__in[15:0] = or_223__out[15:0];
  assign or_225__in0[15:0] = in_450[15:0];
  assign or_225__in1[15:0] = in_451[15:0];
  assign reg_225__in[15:0] = or_225__out[15:0];
  assign or_227__in0[15:0] = in_454[15:0];
  assign or_227__in1[15:0] = in_455[15:0];
  assign reg_227__in[15:0] = or_227__out[15:0];
  assign or_229__in0[15:0] = in_458[15:0];
  assign or_229__in1[15:0] = in_459[15:0];
  assign reg_229__in[15:0] = or_229__out[15:0];
  assign or_23__in0[15:0] = in_46[15:0];
  assign or_23__in1[15:0] = in_47[15:0];
  assign reg_23__in[15:0] = or_23__out[15:0];
  assign or_231__in0[15:0] = in_462[15:0];
  assign or_231__in1[15:0] = in_463[15:0];
  assign reg_231__in[15:0] = or_231__out[15:0];
  assign or_233__in0[15:0] = in_466[15:0];
  assign or_233__in1[15:0] = in_467[15:0];
  assign reg_233__in[15:0] = or_233__out[15:0];
  assign or_235__in0[15:0] = in_470[15:0];
  assign or_235__in1[15:0] = in_471[15:0];
  assign reg_235__in[15:0] = or_235__out[15:0];
  assign or_237__in0[15:0] = in_474[15:0];
  assign or_237__in1[15:0] = in_475[15:0];
  assign reg_237__in[15:0] = or_237__out[15:0];
  assign or_239__in0[15:0] = in_478[15:0];
  assign or_239__in1[15:0] = in_479[15:0];
  assign reg_239__in[15:0] = or_239__out[15:0];
  assign or_241__in0[15:0] = in_482[15:0];
  assign or_241__in1[15:0] = in_483[15:0];
  assign reg_241__in[15:0] = or_241__out[15:0];
  assign or_243__in0[15:0] = in_486[15:0];
  assign or_243__in1[15:0] = in_487[15:0];
  assign reg_243__in[15:0] = or_243__out[15:0];
  assign or_245__in0[15:0] = in_490[15:0];
  assign or_245__in1[15:0] = in_491[15:0];
  assign reg_245__in[15:0] = or_245__out[15:0];
  assign or_247__in0[15:0] = in_494[15:0];
  assign or_247__in1[15:0] = in_495[15:0];
  assign reg_247__in[15:0] = or_247__out[15:0];
  assign or_249__in0[15:0] = in_498[15:0];
  assign or_249__in1[15:0] = in_499[15:0];
  assign reg_249__in[15:0] = or_249__out[15:0];
  assign or_25__in0[15:0] = in_50[15:0];
  assign or_25__in1[15:0] = in_51[15:0];
  assign reg_25__in[15:0] = or_25__out[15:0];
  assign or_251__in0[15:0] = in_502[15:0];
  assign or_251__in1[15:0] = in_503[15:0];
  assign reg_251__in[15:0] = or_251__out[15:0];
  assign or_253__in0[15:0] = in_506[15:0];
  assign or_253__in1[15:0] = in_507[15:0];
  assign reg_253__in[15:0] = or_253__out[15:0];
  assign or_255__in0[15:0] = in_510[15:0];
  assign or_255__in1[15:0] = in_511[15:0];
  assign reg_255__in[15:0] = or_255__out[15:0];
  assign or_257__in0[15:0] = in_514[15:0];
  assign or_257__in1[15:0] = in_515[15:0];
  assign reg_257__in[15:0] = or_257__out[15:0];
  assign or_259__in0[15:0] = in_518[15:0];
  assign or_259__in1[15:0] = in_519[15:0];
  assign reg_259__in[15:0] = or_259__out[15:0];
  assign or_261__in0[15:0] = in_522[15:0];
  assign or_261__in1[15:0] = in_523[15:0];
  assign reg_261__in[15:0] = or_261__out[15:0];
  assign or_263__in0[15:0] = in_526[15:0];
  assign or_263__in1[15:0] = in_527[15:0];
  assign reg_263__in[15:0] = or_263__out[15:0];
  assign or_265__in0[15:0] = in_530[15:0];
  assign or_265__in1[15:0] = in_531[15:0];
  assign reg_265__in[15:0] = or_265__out[15:0];
  assign or_267__in0[15:0] = in_534[15:0];
  assign or_267__in1[15:0] = in_535[15:0];
  assign reg_267__in[15:0] = or_267__out[15:0];
  assign or_269__in0[15:0] = in_538[15:0];
  assign or_269__in1[15:0] = in_539[15:0];
  assign reg_269__in[15:0] = or_269__out[15:0];
  assign or_27__in0[15:0] = in_54[15:0];
  assign or_27__in1[15:0] = in_55[15:0];
  assign reg_27__in[15:0] = or_27__out[15:0];
  assign or_271__in0[15:0] = in_542[15:0];
  assign or_271__in1[15:0] = in_543[15:0];
  assign reg_271__in[15:0] = or_271__out[15:0];
  assign or_273__in0[15:0] = in_546[15:0];
  assign or_273__in1[15:0] = in_547[15:0];
  assign reg_273__in[15:0] = or_273__out[15:0];
  assign or_275__in0[15:0] = in_550[15:0];
  assign or_275__in1[15:0] = in_551[15:0];
  assign reg_275__in[15:0] = or_275__out[15:0];
  assign or_277__in0[15:0] = in_554[15:0];
  assign or_277__in1[15:0] = in_555[15:0];
  assign reg_277__in[15:0] = or_277__out[15:0];
  assign or_279__in0[15:0] = in_558[15:0];
  assign or_279__in1[15:0] = in_559[15:0];
  assign reg_279__in[15:0] = or_279__out[15:0];
  assign or_281__in0[15:0] = in_562[15:0];
  assign or_281__in1[15:0] = in_563[15:0];
  assign reg_281__in[15:0] = or_281__out[15:0];
  assign or_283__in0[15:0] = in_566[15:0];
  assign or_283__in1[15:0] = in_567[15:0];
  assign reg_283__in[15:0] = or_283__out[15:0];
  assign or_285__in0[15:0] = in_570[15:0];
  assign or_285__in1[15:0] = in_571[15:0];
  assign reg_285__in[15:0] = or_285__out[15:0];
  assign or_287__in0[15:0] = in_574[15:0];
  assign or_287__in1[15:0] = in_575[15:0];
  assign reg_287__in[15:0] = or_287__out[15:0];
  assign or_289__in0[15:0] = in_578[15:0];
  assign or_289__in1[15:0] = in_579[15:0];
  assign reg_289__in[15:0] = or_289__out[15:0];
  assign or_29__in0[15:0] = in_58[15:0];
  assign or_29__in1[15:0] = in_59[15:0];
  assign reg_29__in[15:0] = or_29__out[15:0];
  assign or_291__in0[15:0] = in_582[15:0];
  assign or_291__in1[15:0] = in_583[15:0];
  assign reg_291__in[15:0] = or_291__out[15:0];
  assign or_293__in0[15:0] = in_586[15:0];
  assign or_293__in1[15:0] = in_587[15:0];
  assign reg_293__in[15:0] = or_293__out[15:0];
  assign or_295__in0[15:0] = in_590[15:0];
  assign or_295__in1[15:0] = in_591[15:0];
  assign reg_295__in[15:0] = or_295__out[15:0];
  assign or_297__in0[15:0] = in_594[15:0];
  assign or_297__in1[15:0] = in_595[15:0];
  assign reg_297__in[15:0] = or_297__out[15:0];
  assign or_299__in0[15:0] = in_598[15:0];
  assign or_299__in1[15:0] = in_599[15:0];
  assign reg_299__in[15:0] = or_299__out[15:0];
  assign or_3__in0[15:0] = in_6[15:0];
  assign or_3__in1[15:0] = in_7[15:0];
  assign reg_3__in[15:0] = or_3__out[15:0];
  assign or_301__in0[15:0] = in_602[15:0];
  assign or_301__in1[15:0] = in_603[15:0];
  assign reg_301__in[15:0] = or_301__out[15:0];
  assign or_303__in0[15:0] = in_606[15:0];
  assign or_303__in1[15:0] = in_607[15:0];
  assign reg_303__in[15:0] = or_303__out[15:0];
  assign or_305__in0[15:0] = in_610[15:0];
  assign or_305__in1[15:0] = in_611[15:0];
  assign reg_305__in[15:0] = or_305__out[15:0];
  assign or_307__in0[15:0] = in_614[15:0];
  assign or_307__in1[15:0] = in_615[15:0];
  assign reg_307__in[15:0] = or_307__out[15:0];
  assign or_309__in0[15:0] = in_618[15:0];
  assign or_309__in1[15:0] = in_619[15:0];
  assign reg_309__in[15:0] = or_309__out[15:0];
  assign or_31__in0[15:0] = in_62[15:0];
  assign or_31__in1[15:0] = in_63[15:0];
  assign reg_31__in[15:0] = or_31__out[15:0];
  assign or_311__in0[15:0] = in_622[15:0];
  assign or_311__in1[15:0] = in_623[15:0];
  assign reg_311__in[15:0] = or_311__out[15:0];
  assign or_313__in0[15:0] = in_626[15:0];
  assign or_313__in1[15:0] = in_627[15:0];
  assign reg_313__in[15:0] = or_313__out[15:0];
  assign or_315__in0[15:0] = in_630[15:0];
  assign or_315__in1[15:0] = in_631[15:0];
  assign reg_315__in[15:0] = or_315__out[15:0];
  assign or_317__in0[15:0] = in_634[15:0];
  assign or_317__in1[15:0] = in_635[15:0];
  assign reg_317__in[15:0] = or_317__out[15:0];
  assign or_319__in0[15:0] = in_638[15:0];
  assign or_319__in1[15:0] = in_639[15:0];
  assign reg_319__in[15:0] = or_319__out[15:0];
  assign or_321__in0[15:0] = in_642[15:0];
  assign or_321__in1[15:0] = in_643[15:0];
  assign reg_321__in[15:0] = or_321__out[15:0];
  assign or_323__in0[15:0] = in_646[15:0];
  assign or_323__in1[15:0] = in_647[15:0];
  assign reg_323__in[15:0] = or_323__out[15:0];
  assign or_325__in0[15:0] = in_650[15:0];
  assign or_325__in1[15:0] = in_651[15:0];
  assign reg_325__in[15:0] = or_325__out[15:0];
  assign or_327__in0[15:0] = in_654[15:0];
  assign or_327__in1[15:0] = in_655[15:0];
  assign reg_327__in[15:0] = or_327__out[15:0];
  assign or_329__in0[15:0] = in_658[15:0];
  assign or_329__in1[15:0] = in_659[15:0];
  assign reg_329__in[15:0] = or_329__out[15:0];
  assign or_33__in0[15:0] = in_66[15:0];
  assign or_33__in1[15:0] = in_67[15:0];
  assign reg_33__in[15:0] = or_33__out[15:0];
  assign or_331__in0[15:0] = in_662[15:0];
  assign or_331__in1[15:0] = in_663[15:0];
  assign reg_331__in[15:0] = or_331__out[15:0];
  assign or_333__in0[15:0] = in_666[15:0];
  assign or_333__in1[15:0] = in_667[15:0];
  assign reg_333__in[15:0] = or_333__out[15:0];
  assign or_335__in0[15:0] = in_670[15:0];
  assign or_335__in1[15:0] = in_671[15:0];
  assign reg_335__in[15:0] = or_335__out[15:0];
  assign or_337__in0[15:0] = in_674[15:0];
  assign or_337__in1[15:0] = in_675[15:0];
  assign reg_337__in[15:0] = or_337__out[15:0];
  assign or_339__in0[15:0] = in_678[15:0];
  assign or_339__in1[15:0] = in_679[15:0];
  assign reg_339__in[15:0] = or_339__out[15:0];
  assign or_341__in0[15:0] = in_682[15:0];
  assign or_341__in1[15:0] = in_683[15:0];
  assign reg_341__in[15:0] = or_341__out[15:0];
  assign or_343__in0[15:0] = in_686[15:0];
  assign or_343__in1[15:0] = in_687[15:0];
  assign reg_343__in[15:0] = or_343__out[15:0];
  assign or_345__in0[15:0] = in_690[15:0];
  assign or_345__in1[15:0] = in_691[15:0];
  assign reg_345__in[15:0] = or_345__out[15:0];
  assign or_347__in0[15:0] = in_694[15:0];
  assign or_347__in1[15:0] = in_695[15:0];
  assign reg_347__in[15:0] = or_347__out[15:0];
  assign or_349__in0[15:0] = in_698[15:0];
  assign or_349__in1[15:0] = in_699[15:0];
  assign reg_349__in[15:0] = or_349__out[15:0];
  assign or_35__in0[15:0] = in_70[15:0];
  assign or_35__in1[15:0] = in_71[15:0];
  assign reg_35__in[15:0] = or_35__out[15:0];
  assign or_351__in0[15:0] = in_702[15:0];
  assign or_351__in1[15:0] = in_703[15:0];
  assign reg_351__in[15:0] = or_351__out[15:0];
  assign or_353__in0[15:0] = in_706[15:0];
  assign or_353__in1[15:0] = in_707[15:0];
  assign reg_353__in[15:0] = or_353__out[15:0];
  assign or_355__in0[15:0] = in_710[15:0];
  assign or_355__in1[15:0] = in_711[15:0];
  assign reg_355__in[15:0] = or_355__out[15:0];
  assign or_357__in0[15:0] = in_714[15:0];
  assign or_357__in1[15:0] = in_715[15:0];
  assign reg_357__in[15:0] = or_357__out[15:0];
  assign or_359__in0[15:0] = in_718[15:0];
  assign or_359__in1[15:0] = in_719[15:0];
  assign reg_359__in[15:0] = or_359__out[15:0];
  assign or_361__in0[15:0] = in_722[15:0];
  assign or_361__in1[15:0] = in_723[15:0];
  assign reg_361__in[15:0] = or_361__out[15:0];
  assign or_363__in0[15:0] = in_726[15:0];
  assign or_363__in1[15:0] = in_727[15:0];
  assign reg_363__in[15:0] = or_363__out[15:0];
  assign or_365__in0[15:0] = in_730[15:0];
  assign or_365__in1[15:0] = in_731[15:0];
  assign reg_365__in[15:0] = or_365__out[15:0];
  assign or_367__in0[15:0] = in_734[15:0];
  assign or_367__in1[15:0] = in_735[15:0];
  assign reg_367__in[15:0] = or_367__out[15:0];
  assign or_369__in0[15:0] = in_738[15:0];
  assign or_369__in1[15:0] = in_739[15:0];
  assign reg_369__in[15:0] = or_369__out[15:0];
  assign or_37__in0[15:0] = in_74[15:0];
  assign or_37__in1[15:0] = in_75[15:0];
  assign reg_37__in[15:0] = or_37__out[15:0];
  assign or_371__in0[15:0] = in_742[15:0];
  assign or_371__in1[15:0] = in_743[15:0];
  assign reg_371__in[15:0] = or_371__out[15:0];
  assign or_373__in0[15:0] = in_746[15:0];
  assign or_373__in1[15:0] = in_747[15:0];
  assign reg_373__in[15:0] = or_373__out[15:0];
  assign or_375__in0[15:0] = in_750[15:0];
  assign or_375__in1[15:0] = in_751[15:0];
  assign reg_375__in[15:0] = or_375__out[15:0];
  assign or_377__in0[15:0] = in_754[15:0];
  assign or_377__in1[15:0] = in_755[15:0];
  assign reg_377__in[15:0] = or_377__out[15:0];
  assign or_379__in0[15:0] = in_758[15:0];
  assign or_379__in1[15:0] = in_759[15:0];
  assign reg_379__in[15:0] = or_379__out[15:0];
  assign or_381__in0[15:0] = in_762[15:0];
  assign or_381__in1[15:0] = in_763[15:0];
  assign reg_381__in[15:0] = or_381__out[15:0];
  assign or_383__in0[15:0] = in_766[15:0];
  assign or_383__in1[15:0] = in_767[15:0];
  assign reg_383__in[15:0] = or_383__out[15:0];
  assign or_385__in0[15:0] = in_770[15:0];
  assign or_385__in1[15:0] = in_771[15:0];
  assign reg_385__in[15:0] = or_385__out[15:0];
  assign or_387__in0[15:0] = in_774[15:0];
  assign or_387__in1[15:0] = in_775[15:0];
  assign reg_387__in[15:0] = or_387__out[15:0];
  assign or_389__in0[15:0] = in_778[15:0];
  assign or_389__in1[15:0] = in_779[15:0];
  assign reg_389__in[15:0] = or_389__out[15:0];
  assign or_39__in0[15:0] = in_78[15:0];
  assign or_39__in1[15:0] = in_79[15:0];
  assign reg_39__in[15:0] = or_39__out[15:0];
  assign or_391__in0[15:0] = in_782[15:0];
  assign or_391__in1[15:0] = in_783[15:0];
  assign reg_391__in[15:0] = or_391__out[15:0];
  assign or_393__in0[15:0] = in_786[15:0];
  assign or_393__in1[15:0] = in_787[15:0];
  assign reg_393__in[15:0] = or_393__out[15:0];
  assign or_395__in0[15:0] = in_790[15:0];
  assign or_395__in1[15:0] = in_791[15:0];
  assign reg_395__in[15:0] = or_395__out[15:0];
  assign or_397__in0[15:0] = in_794[15:0];
  assign or_397__in1[15:0] = in_795[15:0];
  assign reg_397__in[15:0] = or_397__out[15:0];
  assign or_399__in0[15:0] = in_798[15:0];
  assign or_399__in1[15:0] = in_799[15:0];
  assign reg_399__in[15:0] = or_399__out[15:0];
  assign or_401__in0[15:0] = in_802[15:0];
  assign or_401__in1[15:0] = in_803[15:0];
  assign reg_401__in[15:0] = or_401__out[15:0];
  assign or_403__in0[15:0] = in_806[15:0];
  assign or_403__in1[15:0] = in_807[15:0];
  assign reg_403__in[15:0] = or_403__out[15:0];
  assign or_405__in0[15:0] = in_810[15:0];
  assign or_405__in1[15:0] = in_811[15:0];
  assign reg_405__in[15:0] = or_405__out[15:0];
  assign or_407__in0[15:0] = in_814[15:0];
  assign or_407__in1[15:0] = in_815[15:0];
  assign reg_407__in[15:0] = or_407__out[15:0];
  assign or_409__in0[15:0] = in_818[15:0];
  assign or_409__in1[15:0] = in_819[15:0];
  assign reg_409__in[15:0] = or_409__out[15:0];
  assign or_41__in0[15:0] = in_82[15:0];
  assign or_41__in1[15:0] = in_83[15:0];
  assign reg_41__in[15:0] = or_41__out[15:0];
  assign or_411__in0[15:0] = in_822[15:0];
  assign or_411__in1[15:0] = in_823[15:0];
  assign reg_411__in[15:0] = or_411__out[15:0];
  assign or_413__in0[15:0] = in_826[15:0];
  assign or_413__in1[15:0] = in_827[15:0];
  assign reg_413__in[15:0] = or_413__out[15:0];
  assign or_415__in0[15:0] = in_830[15:0];
  assign or_415__in1[15:0] = in_831[15:0];
  assign reg_415__in[15:0] = or_415__out[15:0];
  assign or_417__in0[15:0] = in_834[15:0];
  assign or_417__in1[15:0] = in_835[15:0];
  assign reg_417__in[15:0] = or_417__out[15:0];
  assign or_419__in0[15:0] = in_838[15:0];
  assign or_419__in1[15:0] = in_839[15:0];
  assign reg_419__in[15:0] = or_419__out[15:0];
  assign or_421__in0[15:0] = in_842[15:0];
  assign or_421__in1[15:0] = in_843[15:0];
  assign reg_421__in[15:0] = or_421__out[15:0];
  assign or_423__in0[15:0] = in_846[15:0];
  assign or_423__in1[15:0] = in_847[15:0];
  assign reg_423__in[15:0] = or_423__out[15:0];
  assign or_425__in0[15:0] = in_850[15:0];
  assign or_425__in1[15:0] = in_851[15:0];
  assign reg_425__in[15:0] = or_425__out[15:0];
  assign or_427__in0[15:0] = in_854[15:0];
  assign or_427__in1[15:0] = in_855[15:0];
  assign reg_427__in[15:0] = or_427__out[15:0];
  assign or_429__in0[15:0] = in_858[15:0];
  assign or_429__in1[15:0] = in_859[15:0];
  assign reg_429__in[15:0] = or_429__out[15:0];
  assign or_43__in0[15:0] = in_86[15:0];
  assign or_43__in1[15:0] = in_87[15:0];
  assign reg_43__in[15:0] = or_43__out[15:0];
  assign or_431__in0[15:0] = in_862[15:0];
  assign or_431__in1[15:0] = in_863[15:0];
  assign reg_431__in[15:0] = or_431__out[15:0];
  assign or_433__in0[15:0] = in_866[15:0];
  assign or_433__in1[15:0] = in_867[15:0];
  assign reg_433__in[15:0] = or_433__out[15:0];
  assign or_435__in0[15:0] = in_870[15:0];
  assign or_435__in1[15:0] = in_871[15:0];
  assign reg_435__in[15:0] = or_435__out[15:0];
  assign or_437__in0[15:0] = in_874[15:0];
  assign or_437__in1[15:0] = in_875[15:0];
  assign reg_437__in[15:0] = or_437__out[15:0];
  assign or_439__in0[15:0] = in_878[15:0];
  assign or_439__in1[15:0] = in_879[15:0];
  assign reg_439__in[15:0] = or_439__out[15:0];
  assign or_441__in0[15:0] = in_882[15:0];
  assign or_441__in1[15:0] = in_883[15:0];
  assign reg_441__in[15:0] = or_441__out[15:0];
  assign or_443__in0[15:0] = in_886[15:0];
  assign or_443__in1[15:0] = in_887[15:0];
  assign reg_443__in[15:0] = or_443__out[15:0];
  assign or_445__in0[15:0] = in_890[15:0];
  assign or_445__in1[15:0] = in_891[15:0];
  assign reg_445__in[15:0] = or_445__out[15:0];
  assign or_447__in0[15:0] = in_894[15:0];
  assign or_447__in1[15:0] = in_895[15:0];
  assign reg_447__in[15:0] = or_447__out[15:0];
  assign or_449__in0[15:0] = in_898[15:0];
  assign or_449__in1[15:0] = in_899[15:0];
  assign reg_449__in[15:0] = or_449__out[15:0];
  assign or_45__in0[15:0] = in_90[15:0];
  assign or_45__in1[15:0] = in_91[15:0];
  assign reg_45__in[15:0] = or_45__out[15:0];
  assign or_451__in0[15:0] = in_902[15:0];
  assign or_451__in1[15:0] = in_903[15:0];
  assign reg_451__in[15:0] = or_451__out[15:0];
  assign or_453__in0[15:0] = in_906[15:0];
  assign or_453__in1[15:0] = in_907[15:0];
  assign reg_453__in[15:0] = or_453__out[15:0];
  assign or_455__in0[15:0] = in_910[15:0];
  assign or_455__in1[15:0] = in_911[15:0];
  assign reg_455__in[15:0] = or_455__out[15:0];
  assign or_457__in0[15:0] = in_914[15:0];
  assign or_457__in1[15:0] = in_915[15:0];
  assign reg_457__in[15:0] = or_457__out[15:0];
  assign or_459__in0[15:0] = in_918[15:0];
  assign or_459__in1[15:0] = in_919[15:0];
  assign reg_459__in[15:0] = or_459__out[15:0];
  assign or_461__in0[15:0] = in_922[15:0];
  assign or_461__in1[15:0] = in_923[15:0];
  assign reg_461__in[15:0] = or_461__out[15:0];
  assign or_463__in0[15:0] = in_926[15:0];
  assign or_463__in1[15:0] = in_927[15:0];
  assign reg_463__in[15:0] = or_463__out[15:0];
  assign or_465__in0[15:0] = in_930[15:0];
  assign or_465__in1[15:0] = in_931[15:0];
  assign reg_465__in[15:0] = or_465__out[15:0];
  assign or_467__in0[15:0] = in_934[15:0];
  assign or_467__in1[15:0] = in_935[15:0];
  assign reg_467__in[15:0] = or_467__out[15:0];
  assign or_469__in0[15:0] = in_938[15:0];
  assign or_469__in1[15:0] = in_939[15:0];
  assign reg_469__in[15:0] = or_469__out[15:0];
  assign or_47__in0[15:0] = in_94[15:0];
  assign or_47__in1[15:0] = in_95[15:0];
  assign reg_47__in[15:0] = or_47__out[15:0];
  assign or_471__in0[15:0] = in_942[15:0];
  assign or_471__in1[15:0] = in_943[15:0];
  assign reg_471__in[15:0] = or_471__out[15:0];
  assign or_473__in0[15:0] = in_946[15:0];
  assign or_473__in1[15:0] = in_947[15:0];
  assign reg_473__in[15:0] = or_473__out[15:0];
  assign or_475__in0[15:0] = in_950[15:0];
  assign or_475__in1[15:0] = in_951[15:0];
  assign reg_475__in[15:0] = or_475__out[15:0];
  assign or_477__in0[15:0] = in_954[15:0];
  assign or_477__in1[15:0] = in_955[15:0];
  assign reg_477__in[15:0] = or_477__out[15:0];
  assign or_479__in0[15:0] = in_958[15:0];
  assign or_479__in1[15:0] = in_959[15:0];
  assign reg_479__in[15:0] = or_479__out[15:0];
  assign or_481__in0[15:0] = in_962[15:0];
  assign or_481__in1[15:0] = in_963[15:0];
  assign reg_481__in[15:0] = or_481__out[15:0];
  assign or_483__in0[15:0] = in_966[15:0];
  assign or_483__in1[15:0] = in_967[15:0];
  assign reg_483__in[15:0] = or_483__out[15:0];
  assign or_485__in0[15:0] = in_970[15:0];
  assign or_485__in1[15:0] = in_971[15:0];
  assign reg_485__in[15:0] = or_485__out[15:0];
  assign or_487__in0[15:0] = in_974[15:0];
  assign or_487__in1[15:0] = in_975[15:0];
  assign reg_487__in[15:0] = or_487__out[15:0];
  assign or_489__in0[15:0] = in_978[15:0];
  assign or_489__in1[15:0] = in_979[15:0];
  assign reg_489__in[15:0] = or_489__out[15:0];
  assign or_49__in0[15:0] = in_98[15:0];
  assign or_49__in1[15:0] = in_99[15:0];
  assign reg_49__in[15:0] = or_49__out[15:0];
  assign or_491__in0[15:0] = in_982[15:0];
  assign or_491__in1[15:0] = in_983[15:0];
  assign reg_491__in[15:0] = or_491__out[15:0];
  assign or_493__in0[15:0] = in_986[15:0];
  assign or_493__in1[15:0] = in_987[15:0];
  assign reg_493__in[15:0] = or_493__out[15:0];
  assign or_495__in0[15:0] = in_990[15:0];
  assign or_495__in1[15:0] = in_991[15:0];
  assign reg_495__in[15:0] = or_495__out[15:0];
  assign or_497__in0[15:0] = in_994[15:0];
  assign or_497__in1[15:0] = in_995[15:0];
  assign reg_497__in[15:0] = or_497__out[15:0];
  assign or_499__in0[15:0] = in_998[15:0];
  assign or_499__in1[15:0] = in_999[15:0];
  assign reg_499__in[15:0] = or_499__out[15:0];
  assign or_5__in0[15:0] = in_10[15:0];
  assign or_5__in1[15:0] = in_11[15:0];
  assign reg_5__in[15:0] = or_5__out[15:0];
  assign or_501__in0[15:0] = in_1002[15:0];
  assign or_501__in1[15:0] = in_1003[15:0];
  assign reg_501__in[15:0] = or_501__out[15:0];
  assign or_503__in0[15:0] = in_1006[15:0];
  assign or_503__in1[15:0] = in_1007[15:0];
  assign reg_503__in[15:0] = or_503__out[15:0];
  assign or_505__in0[15:0] = in_1010[15:0];
  assign or_505__in1[15:0] = in_1011[15:0];
  assign reg_505__in[15:0] = or_505__out[15:0];
  assign or_507__in0[15:0] = in_1014[15:0];
  assign or_507__in1[15:0] = in_1015[15:0];
  assign reg_507__in[15:0] = or_507__out[15:0];
  assign or_509__in0[15:0] = in_1018[15:0];
  assign or_509__in1[15:0] = in_1019[15:0];
  assign reg_509__in[15:0] = or_509__out[15:0];
  assign or_51__in0[15:0] = in_102[15:0];
  assign or_51__in1[15:0] = in_103[15:0];
  assign reg_51__in[15:0] = or_51__out[15:0];
  assign or_511__in0[15:0] = in_1022[15:0];
  assign or_511__in1[15:0] = in_1023[15:0];
  assign reg_511__in[15:0] = or_511__out[15:0];
  assign or_513__in0[15:0] = in_1026[15:0];
  assign or_513__in1[15:0] = in_1027[15:0];
  assign reg_513__in[15:0] = or_513__out[15:0];
  assign or_515__in0[15:0] = in_1030[15:0];
  assign or_515__in1[15:0] = in_1031[15:0];
  assign reg_515__in[15:0] = or_515__out[15:0];
  assign or_517__in0[15:0] = in_1034[15:0];
  assign or_517__in1[15:0] = in_1035[15:0];
  assign reg_517__in[15:0] = or_517__out[15:0];
  assign or_519__in0[15:0] = in_1038[15:0];
  assign or_519__in1[15:0] = in_1039[15:0];
  assign reg_519__in[15:0] = or_519__out[15:0];
  assign or_521__in0[15:0] = in_1042[15:0];
  assign or_521__in1[15:0] = in_1043[15:0];
  assign reg_521__in[15:0] = or_521__out[15:0];
  assign or_523__in0[15:0] = in_1046[15:0];
  assign or_523__in1[15:0] = in_1047[15:0];
  assign reg_523__in[15:0] = or_523__out[15:0];
  assign or_525__in0[15:0] = in_1050[15:0];
  assign or_525__in1[15:0] = in_1051[15:0];
  assign reg_525__in[15:0] = or_525__out[15:0];
  assign or_527__in0[15:0] = in_1054[15:0];
  assign or_527__in1[15:0] = in_1055[15:0];
  assign reg_527__in[15:0] = or_527__out[15:0];
  assign or_529__in0[15:0] = in_1058[15:0];
  assign or_529__in1[15:0] = in_1059[15:0];
  assign reg_529__in[15:0] = or_529__out[15:0];
  assign or_53__in0[15:0] = in_106[15:0];
  assign or_53__in1[15:0] = in_107[15:0];
  assign reg_53__in[15:0] = or_53__out[15:0];
  assign or_531__in0[15:0] = in_1062[15:0];
  assign or_531__in1[15:0] = in_1063[15:0];
  assign reg_531__in[15:0] = or_531__out[15:0];
  assign or_533__in0[15:0] = in_1066[15:0];
  assign or_533__in1[15:0] = in_1067[15:0];
  assign reg_533__in[15:0] = or_533__out[15:0];
  assign or_535__in0[15:0] = in_1070[15:0];
  assign or_535__in1[15:0] = in_1071[15:0];
  assign reg_535__in[15:0] = or_535__out[15:0];
  assign or_537__in0[15:0] = in_1074[15:0];
  assign or_537__in1[15:0] = in_1075[15:0];
  assign reg_537__in[15:0] = or_537__out[15:0];
  assign or_539__in0[15:0] = in_1078[15:0];
  assign or_539__in1[15:0] = in_1079[15:0];
  assign reg_539__in[15:0] = or_539__out[15:0];
  assign or_541__in0[15:0] = in_1082[15:0];
  assign or_541__in1[15:0] = in_1083[15:0];
  assign reg_541__in[15:0] = or_541__out[15:0];
  assign or_543__in0[15:0] = in_1086[15:0];
  assign or_543__in1[15:0] = in_1087[15:0];
  assign reg_543__in[15:0] = or_543__out[15:0];
  assign or_545__in0[15:0] = in_1090[15:0];
  assign or_545__in1[15:0] = in_1091[15:0];
  assign reg_545__in[15:0] = or_545__out[15:0];
  assign or_547__in0[15:0] = in_1094[15:0];
  assign or_547__in1[15:0] = in_1095[15:0];
  assign reg_547__in[15:0] = or_547__out[15:0];
  assign or_549__in0[15:0] = in_1098[15:0];
  assign or_549__in1[15:0] = in_1099[15:0];
  assign reg_549__in[15:0] = or_549__out[15:0];
  assign or_55__in0[15:0] = in_110[15:0];
  assign or_55__in1[15:0] = in_111[15:0];
  assign reg_55__in[15:0] = or_55__out[15:0];
  assign or_551__in0[15:0] = in_1102[15:0];
  assign or_551__in1[15:0] = in_1103[15:0];
  assign reg_551__in[15:0] = or_551__out[15:0];
  assign or_553__in0[15:0] = in_1106[15:0];
  assign or_553__in1[15:0] = in_1107[15:0];
  assign reg_553__in[15:0] = or_553__out[15:0];
  assign or_555__in0[15:0] = in_1110[15:0];
  assign or_555__in1[15:0] = in_1111[15:0];
  assign reg_555__in[15:0] = or_555__out[15:0];
  assign or_557__in0[15:0] = in_1114[15:0];
  assign or_557__in1[15:0] = in_1115[15:0];
  assign reg_557__in[15:0] = or_557__out[15:0];
  assign or_559__in0[15:0] = in_1118[15:0];
  assign or_559__in1[15:0] = in_1119[15:0];
  assign reg_559__in[15:0] = or_559__out[15:0];
  assign or_561__in0[15:0] = in_1122[15:0];
  assign or_561__in1[15:0] = in_1123[15:0];
  assign reg_561__in[15:0] = or_561__out[15:0];
  assign or_563__in0[15:0] = in_1126[15:0];
  assign or_563__in1[15:0] = in_1127[15:0];
  assign reg_563__in[15:0] = or_563__out[15:0];
  assign or_565__in0[15:0] = in_1130[15:0];
  assign or_565__in1[15:0] = in_1131[15:0];
  assign reg_565__in[15:0] = or_565__out[15:0];
  assign or_567__in0[15:0] = in_1134[15:0];
  assign or_567__in1[15:0] = in_1135[15:0];
  assign reg_567__in[15:0] = or_567__out[15:0];
  assign or_569__in0[15:0] = in_1138[15:0];
  assign or_569__in1[15:0] = in_1139[15:0];
  assign reg_569__in[15:0] = or_569__out[15:0];
  assign or_57__in0[15:0] = in_114[15:0];
  assign or_57__in1[15:0] = in_115[15:0];
  assign reg_57__in[15:0] = or_57__out[15:0];
  assign or_571__in0[15:0] = in_1142[15:0];
  assign or_571__in1[15:0] = in_1143[15:0];
  assign reg_571__in[15:0] = or_571__out[15:0];
  assign or_573__in0[15:0] = in_1146[15:0];
  assign or_573__in1[15:0] = in_1147[15:0];
  assign reg_573__in[15:0] = or_573__out[15:0];
  assign or_575__in0[15:0] = in_1150[15:0];
  assign or_575__in1[15:0] = in_1151[15:0];
  assign reg_575__in[15:0] = or_575__out[15:0];
  assign or_577__in0[15:0] = in_1154[15:0];
  assign or_577__in1[15:0] = in_1155[15:0];
  assign reg_577__in[15:0] = or_577__out[15:0];
  assign or_579__in0[15:0] = in_1158[15:0];
  assign or_579__in1[15:0] = in_1159[15:0];
  assign reg_579__in[15:0] = or_579__out[15:0];
  assign or_581__in0[15:0] = in_1162[15:0];
  assign or_581__in1[15:0] = in_1163[15:0];
  assign reg_581__in[15:0] = or_581__out[15:0];
  assign or_583__in0[15:0] = in_1166[15:0];
  assign or_583__in1[15:0] = in_1167[15:0];
  assign reg_583__in[15:0] = or_583__out[15:0];
  assign or_585__in0[15:0] = in_1170[15:0];
  assign or_585__in1[15:0] = in_1171[15:0];
  assign reg_585__in[15:0] = or_585__out[15:0];
  assign or_587__in0[15:0] = in_1174[15:0];
  assign or_587__in1[15:0] = in_1175[15:0];
  assign reg_587__in[15:0] = or_587__out[15:0];
  assign or_589__in0[15:0] = in_1178[15:0];
  assign or_589__in1[15:0] = in_1179[15:0];
  assign reg_589__in[15:0] = or_589__out[15:0];
  assign or_59__in0[15:0] = in_118[15:0];
  assign or_59__in1[15:0] = in_119[15:0];
  assign reg_59__in[15:0] = or_59__out[15:0];
  assign or_591__in0[15:0] = in_1182[15:0];
  assign or_591__in1[15:0] = in_1183[15:0];
  assign reg_591__in[15:0] = or_591__out[15:0];
  assign or_593__in0[15:0] = in_1186[15:0];
  assign or_593__in1[15:0] = in_1187[15:0];
  assign reg_593__in[15:0] = or_593__out[15:0];
  assign or_595__in0[15:0] = in_1190[15:0];
  assign or_595__in1[15:0] = in_1191[15:0];
  assign reg_595__in[15:0] = or_595__out[15:0];
  assign or_597__in0[15:0] = in_1194[15:0];
  assign or_597__in1[15:0] = in_1195[15:0];
  assign reg_597__in[15:0] = or_597__out[15:0];
  assign or_599__in0[15:0] = in_1198[15:0];
  assign or_599__in1[15:0] = in_1199[15:0];
  assign reg_599__in[15:0] = or_599__out[15:0];
  assign or_601__in0[15:0] = in_1202[15:0];
  assign or_601__in1[15:0] = in_1203[15:0];
  assign reg_601__in[15:0] = or_601__out[15:0];
  assign or_603__in0[15:0] = in_1206[15:0];
  assign or_603__in1[15:0] = in_1207[15:0];
  assign reg_603__in[15:0] = or_603__out[15:0];
  assign or_605__in0[15:0] = in_1210[15:0];
  assign or_605__in1[15:0] = in_1211[15:0];
  assign reg_605__in[15:0] = or_605__out[15:0];
  assign or_607__in0[15:0] = in_1214[15:0];
  assign or_607__in1[15:0] = in_1215[15:0];
  assign reg_607__in[15:0] = or_607__out[15:0];
  assign or_609__in0[15:0] = in_1218[15:0];
  assign or_609__in1[15:0] = in_1219[15:0];
  assign reg_609__in[15:0] = or_609__out[15:0];
  assign or_61__in0[15:0] = in_122[15:0];
  assign or_61__in1[15:0] = in_123[15:0];
  assign reg_61__in[15:0] = or_61__out[15:0];
  assign or_611__in0[15:0] = in_1222[15:0];
  assign or_611__in1[15:0] = in_1223[15:0];
  assign reg_611__in[15:0] = or_611__out[15:0];
  assign or_613__in0[15:0] = in_1226[15:0];
  assign or_613__in1[15:0] = in_1227[15:0];
  assign reg_613__in[15:0] = or_613__out[15:0];
  assign or_615__in0[15:0] = in_1230[15:0];
  assign or_615__in1[15:0] = in_1231[15:0];
  assign reg_615__in[15:0] = or_615__out[15:0];
  assign or_617__in0[15:0] = in_1234[15:0];
  assign or_617__in1[15:0] = in_1235[15:0];
  assign reg_617__in[15:0] = or_617__out[15:0];
  assign or_619__in0[15:0] = in_1238[15:0];
  assign or_619__in1[15:0] = in_1239[15:0];
  assign reg_619__in[15:0] = or_619__out[15:0];
  assign or_621__in0[15:0] = in_1242[15:0];
  assign or_621__in1[15:0] = in_1243[15:0];
  assign reg_621__in[15:0] = or_621__out[15:0];
  assign or_623__in0[15:0] = in_1246[15:0];
  assign or_623__in1[15:0] = in_1247[15:0];
  assign reg_623__in[15:0] = or_623__out[15:0];
  assign or_625__in0[15:0] = in_1250[15:0];
  assign or_625__in1[15:0] = in_1251[15:0];
  assign reg_625__in[15:0] = or_625__out[15:0];
  assign or_627__in0[15:0] = in_1254[15:0];
  assign or_627__in1[15:0] = in_1255[15:0];
  assign reg_627__in[15:0] = or_627__out[15:0];
  assign or_629__in0[15:0] = in_1258[15:0];
  assign or_629__in1[15:0] = in_1259[15:0];
  assign reg_629__in[15:0] = or_629__out[15:0];
  assign or_63__in0[15:0] = in_126[15:0];
  assign or_63__in1[15:0] = in_127[15:0];
  assign reg_63__in[15:0] = or_63__out[15:0];
  assign or_631__in0[15:0] = in_1262[15:0];
  assign or_631__in1[15:0] = in_1263[15:0];
  assign reg_631__in[15:0] = or_631__out[15:0];
  assign or_633__in0[15:0] = in_1266[15:0];
  assign or_633__in1[15:0] = in_1267[15:0];
  assign reg_633__in[15:0] = or_633__out[15:0];
  assign or_635__in0[15:0] = in_1270[15:0];
  assign or_635__in1[15:0] = in_1271[15:0];
  assign reg_635__in[15:0] = or_635__out[15:0];
  assign or_637__in0[15:0] = in_1274[15:0];
  assign or_637__in1[15:0] = in_1275[15:0];
  assign reg_637__in[15:0] = or_637__out[15:0];
  assign or_639__in0[15:0] = in_1278[15:0];
  assign or_639__in1[15:0] = in_1279[15:0];
  assign reg_639__in[15:0] = or_639__out[15:0];
  assign or_641__in0[15:0] = in_1282[15:0];
  assign or_641__in1[15:0] = in_1283[15:0];
  assign reg_641__in[15:0] = or_641__out[15:0];
  assign or_643__in0[15:0] = in_1286[15:0];
  assign or_643__in1[15:0] = in_1287[15:0];
  assign reg_643__in[15:0] = or_643__out[15:0];
  assign or_645__in0[15:0] = in_1290[15:0];
  assign or_645__in1[15:0] = in_1291[15:0];
  assign reg_645__in[15:0] = or_645__out[15:0];
  assign or_647__in0[15:0] = in_1294[15:0];
  assign or_647__in1[15:0] = in_1295[15:0];
  assign reg_647__in[15:0] = or_647__out[15:0];
  assign or_649__in0[15:0] = in_1298[15:0];
  assign or_649__in1[15:0] = in_1299[15:0];
  assign reg_649__in[15:0] = or_649__out[15:0];
  assign or_65__in0[15:0] = in_130[15:0];
  assign or_65__in1[15:0] = in_131[15:0];
  assign reg_65__in[15:0] = or_65__out[15:0];
  assign or_651__in0[15:0] = in_1302[15:0];
  assign or_651__in1[15:0] = in_1303[15:0];
  assign reg_651__in[15:0] = or_651__out[15:0];
  assign or_653__in0[15:0] = in_1306[15:0];
  assign or_653__in1[15:0] = in_1307[15:0];
  assign reg_653__in[15:0] = or_653__out[15:0];
  assign or_655__in0[15:0] = in_1310[15:0];
  assign or_655__in1[15:0] = in_1311[15:0];
  assign reg_655__in[15:0] = or_655__out[15:0];
  assign or_657__in0[15:0] = in_1314[15:0];
  assign or_657__in1[15:0] = in_1315[15:0];
  assign reg_657__in[15:0] = or_657__out[15:0];
  assign or_659__in0[15:0] = in_1318[15:0];
  assign or_659__in1[15:0] = in_1319[15:0];
  assign reg_659__in[15:0] = or_659__out[15:0];
  assign or_661__in0[15:0] = in_1322[15:0];
  assign or_661__in1[15:0] = in_1323[15:0];
  assign reg_661__in[15:0] = or_661__out[15:0];
  assign or_663__in0[15:0] = in_1326[15:0];
  assign or_663__in1[15:0] = in_1327[15:0];
  assign reg_663__in[15:0] = or_663__out[15:0];
  assign or_665__in0[15:0] = in_1330[15:0];
  assign or_665__in1[15:0] = in_1331[15:0];
  assign reg_665__in[15:0] = or_665__out[15:0];
  assign or_667__in0[15:0] = in_1334[15:0];
  assign or_667__in1[15:0] = in_1335[15:0];
  assign reg_667__in[15:0] = or_667__out[15:0];
  assign or_669__in0[15:0] = in_1338[15:0];
  assign or_669__in1[15:0] = in_1339[15:0];
  assign reg_669__in[15:0] = or_669__out[15:0];
  assign or_67__in0[15:0] = in_134[15:0];
  assign or_67__in1[15:0] = in_135[15:0];
  assign reg_67__in[15:0] = or_67__out[15:0];
  assign or_671__in0[15:0] = in_1342[15:0];
  assign or_671__in1[15:0] = in_1343[15:0];
  assign reg_671__in[15:0] = or_671__out[15:0];
  assign or_673__in0[15:0] = in_1346[15:0];
  assign or_673__in1[15:0] = in_1347[15:0];
  assign reg_673__in[15:0] = or_673__out[15:0];
  assign or_675__in0[15:0] = in_1350[15:0];
  assign or_675__in1[15:0] = in_1351[15:0];
  assign reg_675__in[15:0] = or_675__out[15:0];
  assign or_677__in0[15:0] = in_1354[15:0];
  assign or_677__in1[15:0] = in_1355[15:0];
  assign reg_677__in[15:0] = or_677__out[15:0];
  assign or_679__in0[15:0] = in_1358[15:0];
  assign or_679__in1[15:0] = in_1359[15:0];
  assign reg_679__in[15:0] = or_679__out[15:0];
  assign or_681__in0[15:0] = in_1362[15:0];
  assign or_681__in1[15:0] = in_1363[15:0];
  assign reg_681__in[15:0] = or_681__out[15:0];
  assign or_683__in0[15:0] = in_1366[15:0];
  assign or_683__in1[15:0] = in_1367[15:0];
  assign reg_683__in[15:0] = or_683__out[15:0];
  assign or_685__in0[15:0] = in_1370[15:0];
  assign or_685__in1[15:0] = in_1371[15:0];
  assign reg_685__in[15:0] = or_685__out[15:0];
  assign or_687__in0[15:0] = in_1374[15:0];
  assign or_687__in1[15:0] = in_1375[15:0];
  assign reg_687__in[15:0] = or_687__out[15:0];
  assign or_689__in0[15:0] = in_1378[15:0];
  assign or_689__in1[15:0] = in_1379[15:0];
  assign reg_689__in[15:0] = or_689__out[15:0];
  assign or_69__in0[15:0] = in_138[15:0];
  assign or_69__in1[15:0] = in_139[15:0];
  assign reg_69__in[15:0] = or_69__out[15:0];
  assign or_691__in0[15:0] = in_1382[15:0];
  assign or_691__in1[15:0] = in_1383[15:0];
  assign reg_691__in[15:0] = or_691__out[15:0];
  assign or_693__in0[15:0] = in_1386[15:0];
  assign or_693__in1[15:0] = in_1387[15:0];
  assign reg_693__in[15:0] = or_693__out[15:0];
  assign or_695__in0[15:0] = in_1390[15:0];
  assign or_695__in1[15:0] = in_1391[15:0];
  assign reg_695__in[15:0] = or_695__out[15:0];
  assign or_697__in0[15:0] = in_1394[15:0];
  assign or_697__in1[15:0] = in_1395[15:0];
  assign reg_697__in[15:0] = or_697__out[15:0];
  assign or_699__in0[15:0] = in_1398[15:0];
  assign or_699__in1[15:0] = in_1399[15:0];
  assign reg_699__in[15:0] = or_699__out[15:0];
  assign or_7__in0[15:0] = in_14[15:0];
  assign or_7__in1[15:0] = in_15[15:0];
  assign reg_7__in[15:0] = or_7__out[15:0];
  assign or_701__in0[15:0] = in_1402[15:0];
  assign or_701__in1[15:0] = in_1403[15:0];
  assign reg_701__in[15:0] = or_701__out[15:0];
  assign or_703__in0[15:0] = in_1406[15:0];
  assign or_703__in1[15:0] = in_1407[15:0];
  assign reg_703__in[15:0] = or_703__out[15:0];
  assign or_705__in0[15:0] = in_1410[15:0];
  assign or_705__in1[15:0] = in_1411[15:0];
  assign reg_705__in[15:0] = or_705__out[15:0];
  assign or_707__in0[15:0] = in_1414[15:0];
  assign or_707__in1[15:0] = in_1415[15:0];
  assign reg_707__in[15:0] = or_707__out[15:0];
  assign or_709__in0[15:0] = in_1418[15:0];
  assign or_709__in1[15:0] = in_1419[15:0];
  assign reg_709__in[15:0] = or_709__out[15:0];
  assign or_71__in0[15:0] = in_142[15:0];
  assign or_71__in1[15:0] = in_143[15:0];
  assign reg_71__in[15:0] = or_71__out[15:0];
  assign or_711__in0[15:0] = in_1422[15:0];
  assign or_711__in1[15:0] = in_1423[15:0];
  assign reg_711__in[15:0] = or_711__out[15:0];
  assign or_713__in0[15:0] = in_1426[15:0];
  assign or_713__in1[15:0] = in_1427[15:0];
  assign reg_713__in[15:0] = or_713__out[15:0];
  assign or_715__in0[15:0] = in_1430[15:0];
  assign or_715__in1[15:0] = in_1431[15:0];
  assign reg_715__in[15:0] = or_715__out[15:0];
  assign or_717__in0[15:0] = in_1434[15:0];
  assign or_717__in1[15:0] = in_1435[15:0];
  assign reg_717__in[15:0] = or_717__out[15:0];
  assign or_719__in0[15:0] = in_1438[15:0];
  assign or_719__in1[15:0] = in_1439[15:0];
  assign reg_719__in[15:0] = or_719__out[15:0];
  assign or_721__in0[15:0] = in_1442[15:0];
  assign or_721__in1[15:0] = in_1443[15:0];
  assign reg_721__in[15:0] = or_721__out[15:0];
  assign or_723__in0[15:0] = in_1446[15:0];
  assign or_723__in1[15:0] = in_1447[15:0];
  assign reg_723__in[15:0] = or_723__out[15:0];
  assign or_725__in0[15:0] = in_1450[15:0];
  assign or_725__in1[15:0] = in_1451[15:0];
  assign reg_725__in[15:0] = or_725__out[15:0];
  assign or_727__in0[15:0] = in_1454[15:0];
  assign or_727__in1[15:0] = in_1455[15:0];
  assign reg_727__in[15:0] = or_727__out[15:0];
  assign or_729__in0[15:0] = in_1458[15:0];
  assign or_729__in1[15:0] = in_1459[15:0];
  assign reg_729__in[15:0] = or_729__out[15:0];
  assign or_73__in0[15:0] = in_146[15:0];
  assign or_73__in1[15:0] = in_147[15:0];
  assign reg_73__in[15:0] = or_73__out[15:0];
  assign or_731__in0[15:0] = in_1462[15:0];
  assign or_731__in1[15:0] = in_1463[15:0];
  assign reg_731__in[15:0] = or_731__out[15:0];
  assign or_733__in0[15:0] = in_1466[15:0];
  assign or_733__in1[15:0] = in_1467[15:0];
  assign reg_733__in[15:0] = or_733__out[15:0];
  assign or_735__in0[15:0] = in_1470[15:0];
  assign or_735__in1[15:0] = in_1471[15:0];
  assign reg_735__in[15:0] = or_735__out[15:0];
  assign or_737__in0[15:0] = in_1474[15:0];
  assign or_737__in1[15:0] = in_1475[15:0];
  assign reg_737__in[15:0] = or_737__out[15:0];
  assign or_739__in0[15:0] = in_1478[15:0];
  assign or_739__in1[15:0] = in_1479[15:0];
  assign reg_739__in[15:0] = or_739__out[15:0];
  assign or_741__in0[15:0] = in_1482[15:0];
  assign or_741__in1[15:0] = in_1483[15:0];
  assign reg_741__in[15:0] = or_741__out[15:0];
  assign or_743__in0[15:0] = in_1486[15:0];
  assign or_743__in1[15:0] = in_1487[15:0];
  assign reg_743__in[15:0] = or_743__out[15:0];
  assign or_745__in0[15:0] = in_1490[15:0];
  assign or_745__in1[15:0] = in_1491[15:0];
  assign reg_745__in[15:0] = or_745__out[15:0];
  assign or_747__in0[15:0] = in_1494[15:0];
  assign or_747__in1[15:0] = in_1495[15:0];
  assign reg_747__in[15:0] = or_747__out[15:0];
  assign or_749__in0[15:0] = in_1498[15:0];
  assign or_749__in1[15:0] = in_1499[15:0];
  assign reg_749__in[15:0] = or_749__out[15:0];
  assign or_75__in0[15:0] = in_150[15:0];
  assign or_75__in1[15:0] = in_151[15:0];
  assign reg_75__in[15:0] = or_75__out[15:0];
  assign or_751__in0[15:0] = in_1502[15:0];
  assign or_751__in1[15:0] = in_1503[15:0];
  assign reg_751__in[15:0] = or_751__out[15:0];
  assign or_753__in0[15:0] = in_1506[15:0];
  assign or_753__in1[15:0] = in_1507[15:0];
  assign reg_753__in[15:0] = or_753__out[15:0];
  assign or_755__in0[15:0] = in_1510[15:0];
  assign or_755__in1[15:0] = in_1511[15:0];
  assign reg_755__in[15:0] = or_755__out[15:0];
  assign or_757__in0[15:0] = in_1514[15:0];
  assign or_757__in1[15:0] = in_1515[15:0];
  assign reg_757__in[15:0] = or_757__out[15:0];
  assign or_759__in0[15:0] = in_1518[15:0];
  assign or_759__in1[15:0] = in_1519[15:0];
  assign reg_759__in[15:0] = or_759__out[15:0];
  assign or_761__in0[15:0] = in_1522[15:0];
  assign or_761__in1[15:0] = in_1523[15:0];
  assign reg_761__in[15:0] = or_761__out[15:0];
  assign or_763__in0[15:0] = in_1526[15:0];
  assign or_763__in1[15:0] = in_1527[15:0];
  assign reg_763__in[15:0] = or_763__out[15:0];
  assign or_765__in0[15:0] = in_1530[15:0];
  assign or_765__in1[15:0] = in_1531[15:0];
  assign reg_765__in[15:0] = or_765__out[15:0];
  assign or_767__in0[15:0] = in_1534[15:0];
  assign or_767__in1[15:0] = in_1535[15:0];
  assign reg_767__in[15:0] = or_767__out[15:0];
  assign or_769__in0[15:0] = in_1538[15:0];
  assign or_769__in1[15:0] = in_1539[15:0];
  assign reg_769__in[15:0] = or_769__out[15:0];
  assign or_77__in0[15:0] = in_154[15:0];
  assign or_77__in1[15:0] = in_155[15:0];
  assign reg_77__in[15:0] = or_77__out[15:0];
  assign or_771__in0[15:0] = in_1542[15:0];
  assign or_771__in1[15:0] = in_1543[15:0];
  assign reg_771__in[15:0] = or_771__out[15:0];
  assign or_773__in0[15:0] = in_1546[15:0];
  assign or_773__in1[15:0] = in_1547[15:0];
  assign reg_773__in[15:0] = or_773__out[15:0];
  assign or_775__in0[15:0] = in_1550[15:0];
  assign or_775__in1[15:0] = in_1551[15:0];
  assign reg_775__in[15:0] = or_775__out[15:0];
  assign or_777__in0[15:0] = in_1554[15:0];
  assign or_777__in1[15:0] = in_1555[15:0];
  assign reg_777__in[15:0] = or_777__out[15:0];
  assign or_779__in0[15:0] = in_1558[15:0];
  assign or_779__in1[15:0] = in_1559[15:0];
  assign reg_779__in[15:0] = or_779__out[15:0];
  assign or_781__in0[15:0] = in_1562[15:0];
  assign or_781__in1[15:0] = in_1563[15:0];
  assign reg_781__in[15:0] = or_781__out[15:0];
  assign or_783__in0[15:0] = in_1566[15:0];
  assign or_783__in1[15:0] = in_1567[15:0];
  assign reg_783__in[15:0] = or_783__out[15:0];
  assign or_785__in0[15:0] = in_1570[15:0];
  assign or_785__in1[15:0] = in_1571[15:0];
  assign reg_785__in[15:0] = or_785__out[15:0];
  assign or_787__in0[15:0] = in_1574[15:0];
  assign or_787__in1[15:0] = in_1575[15:0];
  assign reg_787__in[15:0] = or_787__out[15:0];
  assign or_789__in0[15:0] = in_1578[15:0];
  assign or_789__in1[15:0] = in_1579[15:0];
  assign reg_789__in[15:0] = or_789__out[15:0];
  assign or_79__in0[15:0] = in_158[15:0];
  assign or_79__in1[15:0] = in_159[15:0];
  assign reg_79__in[15:0] = or_79__out[15:0];
  assign or_791__in0[15:0] = in_1582[15:0];
  assign or_791__in1[15:0] = in_1583[15:0];
  assign reg_791__in[15:0] = or_791__out[15:0];
  assign or_793__in0[15:0] = in_1586[15:0];
  assign or_793__in1[15:0] = in_1587[15:0];
  assign reg_793__in[15:0] = or_793__out[15:0];
  assign or_795__in0[15:0] = in_1590[15:0];
  assign or_795__in1[15:0] = in_1591[15:0];
  assign reg_795__in[15:0] = or_795__out[15:0];
  assign or_797__in0[15:0] = in_1594[15:0];
  assign or_797__in1[15:0] = in_1595[15:0];
  assign reg_797__in[15:0] = or_797__out[15:0];
  assign or_799__in0[15:0] = in_1598[15:0];
  assign or_799__in1[15:0] = in_1599[15:0];
  assign reg_799__in[15:0] = or_799__out[15:0];
  assign or_801__in0[15:0] = in_1602[15:0];
  assign or_801__in1[15:0] = in_1603[15:0];
  assign reg_801__in[15:0] = or_801__out[15:0];
  assign or_803__in0[15:0] = in_1606[15:0];
  assign or_803__in1[15:0] = in_1607[15:0];
  assign reg_803__in[15:0] = or_803__out[15:0];
  assign or_805__in0[15:0] = in_1610[15:0];
  assign or_805__in1[15:0] = in_1611[15:0];
  assign reg_805__in[15:0] = or_805__out[15:0];
  assign or_807__in0[15:0] = in_1614[15:0];
  assign or_807__in1[15:0] = in_1615[15:0];
  assign reg_807__in[15:0] = or_807__out[15:0];
  assign or_809__in0[15:0] = in_1618[15:0];
  assign or_809__in1[15:0] = in_1619[15:0];
  assign reg_809__in[15:0] = or_809__out[15:0];
  assign or_81__in0[15:0] = in_162[15:0];
  assign or_81__in1[15:0] = in_163[15:0];
  assign reg_81__in[15:0] = or_81__out[15:0];
  assign or_811__in0[15:0] = in_1622[15:0];
  assign or_811__in1[15:0] = in_1623[15:0];
  assign reg_811__in[15:0] = or_811__out[15:0];
  assign or_813__in0[15:0] = in_1626[15:0];
  assign or_813__in1[15:0] = in_1627[15:0];
  assign reg_813__in[15:0] = or_813__out[15:0];
  assign or_815__in0[15:0] = in_1630[15:0];
  assign or_815__in1[15:0] = in_1631[15:0];
  assign reg_815__in[15:0] = or_815__out[15:0];
  assign or_817__in0[15:0] = in_1634[15:0];
  assign or_817__in1[15:0] = in_1635[15:0];
  assign reg_817__in[15:0] = or_817__out[15:0];
  assign or_819__in0[15:0] = in_1638[15:0];
  assign or_819__in1[15:0] = in_1639[15:0];
  assign reg_819__in[15:0] = or_819__out[15:0];
  assign or_821__in0[15:0] = in_1642[15:0];
  assign or_821__in1[15:0] = in_1643[15:0];
  assign reg_821__in[15:0] = or_821__out[15:0];
  assign or_823__in0[15:0] = in_1646[15:0];
  assign or_823__in1[15:0] = in_1647[15:0];
  assign reg_823__in[15:0] = or_823__out[15:0];
  assign or_825__in0[15:0] = in_1650[15:0];
  assign or_825__in1[15:0] = in_1651[15:0];
  assign reg_825__in[15:0] = or_825__out[15:0];
  assign or_827__in0[15:0] = in_1654[15:0];
  assign or_827__in1[15:0] = in_1655[15:0];
  assign reg_827__in[15:0] = or_827__out[15:0];
  assign or_829__in0[15:0] = in_1658[15:0];
  assign or_829__in1[15:0] = in_1659[15:0];
  assign reg_829__in[15:0] = or_829__out[15:0];
  assign or_83__in0[15:0] = in_166[15:0];
  assign or_83__in1[15:0] = in_167[15:0];
  assign reg_83__in[15:0] = or_83__out[15:0];
  assign or_831__in0[15:0] = in_1662[15:0];
  assign or_831__in1[15:0] = in_1663[15:0];
  assign reg_831__in[15:0] = or_831__out[15:0];
  assign or_833__in0[15:0] = in_1666[15:0];
  assign or_833__in1[15:0] = in_1667[15:0];
  assign reg_833__in[15:0] = or_833__out[15:0];
  assign or_835__in0[15:0] = in_1670[15:0];
  assign or_835__in1[15:0] = in_1671[15:0];
  assign reg_835__in[15:0] = or_835__out[15:0];
  assign or_837__in0[15:0] = in_1674[15:0];
  assign or_837__in1[15:0] = in_1675[15:0];
  assign reg_837__in[15:0] = or_837__out[15:0];
  assign or_839__in0[15:0] = in_1678[15:0];
  assign or_839__in1[15:0] = in_1679[15:0];
  assign reg_839__in[15:0] = or_839__out[15:0];
  assign or_841__in0[15:0] = in_1682[15:0];
  assign or_841__in1[15:0] = in_1683[15:0];
  assign reg_841__in[15:0] = or_841__out[15:0];
  assign or_843__in0[15:0] = in_1686[15:0];
  assign or_843__in1[15:0] = in_1687[15:0];
  assign reg_843__in[15:0] = or_843__out[15:0];
  assign or_845__in0[15:0] = in_1690[15:0];
  assign or_845__in1[15:0] = in_1691[15:0];
  assign reg_845__in[15:0] = or_845__out[15:0];
  assign or_847__in0[15:0] = in_1694[15:0];
  assign or_847__in1[15:0] = in_1695[15:0];
  assign reg_847__in[15:0] = or_847__out[15:0];
  assign or_849__in0[15:0] = in_1698[15:0];
  assign or_849__in1[15:0] = in_1699[15:0];
  assign reg_849__in[15:0] = or_849__out[15:0];
  assign or_85__in0[15:0] = in_170[15:0];
  assign or_85__in1[15:0] = in_171[15:0];
  assign reg_85__in[15:0] = or_85__out[15:0];
  assign or_851__in0[15:0] = in_1702[15:0];
  assign or_851__in1[15:0] = in_1703[15:0];
  assign reg_851__in[15:0] = or_851__out[15:0];
  assign or_853__in0[15:0] = in_1706[15:0];
  assign or_853__in1[15:0] = in_1707[15:0];
  assign reg_853__in[15:0] = or_853__out[15:0];
  assign or_855__in0[15:0] = in_1710[15:0];
  assign or_855__in1[15:0] = in_1711[15:0];
  assign reg_855__in[15:0] = or_855__out[15:0];
  assign or_857__in0[15:0] = in_1714[15:0];
  assign or_857__in1[15:0] = in_1715[15:0];
  assign reg_857__in[15:0] = or_857__out[15:0];
  assign or_859__in0[15:0] = in_1718[15:0];
  assign or_859__in1[15:0] = in_1719[15:0];
  assign reg_859__in[15:0] = or_859__out[15:0];
  assign or_861__in0[15:0] = in_1722[15:0];
  assign or_861__in1[15:0] = in_1723[15:0];
  assign reg_861__in[15:0] = or_861__out[15:0];
  assign or_863__in0[15:0] = in_1726[15:0];
  assign or_863__in1[15:0] = in_1727[15:0];
  assign reg_863__in[15:0] = or_863__out[15:0];
  assign or_865__in0[15:0] = in_1730[15:0];
  assign or_865__in1[15:0] = in_1731[15:0];
  assign reg_865__in[15:0] = or_865__out[15:0];
  assign or_867__in0[15:0] = in_1734[15:0];
  assign or_867__in1[15:0] = in_1735[15:0];
  assign reg_867__in[15:0] = or_867__out[15:0];
  assign or_869__in0[15:0] = in_1738[15:0];
  assign or_869__in1[15:0] = in_1739[15:0];
  assign reg_869__in[15:0] = or_869__out[15:0];
  assign or_87__in0[15:0] = in_174[15:0];
  assign or_87__in1[15:0] = in_175[15:0];
  assign reg_87__in[15:0] = or_87__out[15:0];
  assign or_871__in0[15:0] = in_1742[15:0];
  assign or_871__in1[15:0] = in_1743[15:0];
  assign reg_871__in[15:0] = or_871__out[15:0];
  assign or_873__in0[15:0] = in_1746[15:0];
  assign or_873__in1[15:0] = in_1747[15:0];
  assign reg_873__in[15:0] = or_873__out[15:0];
  assign or_875__in0[15:0] = in_1750[15:0];
  assign or_875__in1[15:0] = in_1751[15:0];
  assign reg_875__in[15:0] = or_875__out[15:0];
  assign or_877__in0[15:0] = in_1754[15:0];
  assign or_877__in1[15:0] = in_1755[15:0];
  assign reg_877__in[15:0] = or_877__out[15:0];
  assign or_879__in0[15:0] = in_1758[15:0];
  assign or_879__in1[15:0] = in_1759[15:0];
  assign reg_879__in[15:0] = or_879__out[15:0];
  assign or_881__in0[15:0] = in_1762[15:0];
  assign or_881__in1[15:0] = in_1763[15:0];
  assign reg_881__in[15:0] = or_881__out[15:0];
  assign or_883__in0[15:0] = in_1766[15:0];
  assign or_883__in1[15:0] = in_1767[15:0];
  assign reg_883__in[15:0] = or_883__out[15:0];
  assign or_885__in0[15:0] = in_1770[15:0];
  assign or_885__in1[15:0] = in_1771[15:0];
  assign reg_885__in[15:0] = or_885__out[15:0];
  assign or_887__in0[15:0] = in_1774[15:0];
  assign or_887__in1[15:0] = in_1775[15:0];
  assign reg_887__in[15:0] = or_887__out[15:0];
  assign or_889__in0[15:0] = in_1778[15:0];
  assign or_889__in1[15:0] = in_1779[15:0];
  assign reg_889__in[15:0] = or_889__out[15:0];
  assign or_89__in0[15:0] = in_178[15:0];
  assign or_89__in1[15:0] = in_179[15:0];
  assign reg_89__in[15:0] = or_89__out[15:0];
  assign or_891__in0[15:0] = in_1782[15:0];
  assign or_891__in1[15:0] = in_1783[15:0];
  assign reg_891__in[15:0] = or_891__out[15:0];
  assign or_893__in0[15:0] = in_1786[15:0];
  assign or_893__in1[15:0] = in_1787[15:0];
  assign reg_893__in[15:0] = or_893__out[15:0];
  assign or_895__in0[15:0] = in_1790[15:0];
  assign or_895__in1[15:0] = in_1791[15:0];
  assign reg_895__in[15:0] = or_895__out[15:0];
  assign or_897__in0[15:0] = in_1794[15:0];
  assign or_897__in1[15:0] = in_1795[15:0];
  assign reg_897__in[15:0] = or_897__out[15:0];
  assign or_899__in0[15:0] = in_1798[15:0];
  assign or_899__in1[15:0] = in_1799[15:0];
  assign reg_899__in[15:0] = or_899__out[15:0];
  assign or_9__in0[15:0] = in_18[15:0];
  assign or_9__in1[15:0] = in_19[15:0];
  assign reg_9__in[15:0] = or_9__out[15:0];
  assign or_901__in0[15:0] = in_1802[15:0];
  assign or_901__in1[15:0] = in_1803[15:0];
  assign reg_901__in[15:0] = or_901__out[15:0];
  assign or_903__in0[15:0] = in_1806[15:0];
  assign or_903__in1[15:0] = in_1807[15:0];
  assign reg_903__in[15:0] = or_903__out[15:0];
  assign or_905__in0[15:0] = in_1810[15:0];
  assign or_905__in1[15:0] = in_1811[15:0];
  assign reg_905__in[15:0] = or_905__out[15:0];
  assign or_907__in0[15:0] = in_1814[15:0];
  assign or_907__in1[15:0] = in_1815[15:0];
  assign reg_907__in[15:0] = or_907__out[15:0];
  assign or_909__in0[15:0] = in_1818[15:0];
  assign or_909__in1[15:0] = in_1819[15:0];
  assign reg_909__in[15:0] = or_909__out[15:0];
  assign or_91__in0[15:0] = in_182[15:0];
  assign or_91__in1[15:0] = in_183[15:0];
  assign reg_91__in[15:0] = or_91__out[15:0];
  assign or_911__in0[15:0] = in_1822[15:0];
  assign or_911__in1[15:0] = in_1823[15:0];
  assign reg_911__in[15:0] = or_911__out[15:0];
  assign or_913__in0[15:0] = in_1826[15:0];
  assign or_913__in1[15:0] = in_1827[15:0];
  assign reg_913__in[15:0] = or_913__out[15:0];
  assign or_915__in0[15:0] = in_1830[15:0];
  assign or_915__in1[15:0] = in_1831[15:0];
  assign reg_915__in[15:0] = or_915__out[15:0];
  assign or_917__in0[15:0] = in_1834[15:0];
  assign or_917__in1[15:0] = in_1835[15:0];
  assign reg_917__in[15:0] = or_917__out[15:0];
  assign or_919__in0[15:0] = in_1838[15:0];
  assign or_919__in1[15:0] = in_1839[15:0];
  assign reg_919__in[15:0] = or_919__out[15:0];
  assign or_921__in0[15:0] = in_1842[15:0];
  assign or_921__in1[15:0] = in_1843[15:0];
  assign reg_921__in[15:0] = or_921__out[15:0];
  assign or_923__in0[15:0] = in_1846[15:0];
  assign or_923__in1[15:0] = in_1847[15:0];
  assign reg_923__in[15:0] = or_923__out[15:0];
  assign or_925__in0[15:0] = in_1850[15:0];
  assign or_925__in1[15:0] = in_1851[15:0];
  assign reg_925__in[15:0] = or_925__out[15:0];
  assign or_927__in0[15:0] = in_1854[15:0];
  assign or_927__in1[15:0] = in_1855[15:0];
  assign reg_927__in[15:0] = or_927__out[15:0];
  assign or_929__in0[15:0] = in_1858[15:0];
  assign or_929__in1[15:0] = in_1859[15:0];
  assign reg_929__in[15:0] = or_929__out[15:0];
  assign or_93__in0[15:0] = in_186[15:0];
  assign or_93__in1[15:0] = in_187[15:0];
  assign reg_93__in[15:0] = or_93__out[15:0];
  assign or_931__in0[15:0] = in_1862[15:0];
  assign or_931__in1[15:0] = in_1863[15:0];
  assign reg_931__in[15:0] = or_931__out[15:0];
  assign or_933__in0[15:0] = in_1866[15:0];
  assign or_933__in1[15:0] = in_1867[15:0];
  assign reg_933__in[15:0] = or_933__out[15:0];
  assign or_935__in0[15:0] = in_1870[15:0];
  assign or_935__in1[15:0] = in_1871[15:0];
  assign reg_935__in[15:0] = or_935__out[15:0];
  assign or_937__in0[15:0] = in_1874[15:0];
  assign or_937__in1[15:0] = in_1875[15:0];
  assign reg_937__in[15:0] = or_937__out[15:0];
  assign or_939__in0[15:0] = in_1878[15:0];
  assign or_939__in1[15:0] = in_1879[15:0];
  assign reg_939__in[15:0] = or_939__out[15:0];
  assign or_941__in0[15:0] = in_1882[15:0];
  assign or_941__in1[15:0] = in_1883[15:0];
  assign reg_941__in[15:0] = or_941__out[15:0];
  assign or_943__in0[15:0] = in_1886[15:0];
  assign or_943__in1[15:0] = in_1887[15:0];
  assign reg_943__in[15:0] = or_943__out[15:0];
  assign or_945__in0[15:0] = in_1890[15:0];
  assign or_945__in1[15:0] = in_1891[15:0];
  assign reg_945__in[15:0] = or_945__out[15:0];
  assign or_947__in0[15:0] = in_1894[15:0];
  assign or_947__in1[15:0] = in_1895[15:0];
  assign reg_947__in[15:0] = or_947__out[15:0];
  assign or_949__in0[15:0] = in_1898[15:0];
  assign or_949__in1[15:0] = in_1899[15:0];
  assign reg_949__in[15:0] = or_949__out[15:0];
  assign or_95__in0[15:0] = in_190[15:0];
  assign or_95__in1[15:0] = in_191[15:0];
  assign reg_95__in[15:0] = or_95__out[15:0];
  assign or_951__in0[15:0] = in_1902[15:0];
  assign or_951__in1[15:0] = in_1903[15:0];
  assign reg_951__in[15:0] = or_951__out[15:0];
  assign or_953__in0[15:0] = in_1906[15:0];
  assign or_953__in1[15:0] = in_1907[15:0];
  assign reg_953__in[15:0] = or_953__out[15:0];
  assign or_955__in0[15:0] = in_1910[15:0];
  assign or_955__in1[15:0] = in_1911[15:0];
  assign reg_955__in[15:0] = or_955__out[15:0];
  assign or_957__in0[15:0] = in_1914[15:0];
  assign or_957__in1[15:0] = in_1915[15:0];
  assign reg_957__in[15:0] = or_957__out[15:0];
  assign or_959__in0[15:0] = in_1918[15:0];
  assign or_959__in1[15:0] = in_1919[15:0];
  assign reg_959__in[15:0] = or_959__out[15:0];
  assign or_961__in0[15:0] = in_1922[15:0];
  assign or_961__in1[15:0] = in_1923[15:0];
  assign reg_961__in[15:0] = or_961__out[15:0];
  assign or_963__in0[15:0] = in_1926[15:0];
  assign or_963__in1[15:0] = in_1927[15:0];
  assign reg_963__in[15:0] = or_963__out[15:0];
  assign or_965__in0[15:0] = in_1930[15:0];
  assign or_965__in1[15:0] = in_1931[15:0];
  assign reg_965__in[15:0] = or_965__out[15:0];
  assign or_967__in0[15:0] = in_1934[15:0];
  assign or_967__in1[15:0] = in_1935[15:0];
  assign reg_967__in[15:0] = or_967__out[15:0];
  assign or_969__in0[15:0] = in_1938[15:0];
  assign or_969__in1[15:0] = in_1939[15:0];
  assign reg_969__in[15:0] = or_969__out[15:0];
  assign or_97__in0[15:0] = in_194[15:0];
  assign or_97__in1[15:0] = in_195[15:0];
  assign reg_97__in[15:0] = or_97__out[15:0];
  assign or_971__in0[15:0] = in_1942[15:0];
  assign or_971__in1[15:0] = in_1943[15:0];
  assign reg_971__in[15:0] = or_971__out[15:0];
  assign or_973__in0[15:0] = in_1946[15:0];
  assign or_973__in1[15:0] = in_1947[15:0];
  assign reg_973__in[15:0] = or_973__out[15:0];
  assign or_975__in0[15:0] = in_1950[15:0];
  assign or_975__in1[15:0] = in_1951[15:0];
  assign reg_975__in[15:0] = or_975__out[15:0];
  assign or_977__in0[15:0] = in_1954[15:0];
  assign or_977__in1[15:0] = in_1955[15:0];
  assign reg_977__in[15:0] = or_977__out[15:0];
  assign or_979__in0[15:0] = in_1958[15:0];
  assign or_979__in1[15:0] = in_1959[15:0];
  assign reg_979__in[15:0] = or_979__out[15:0];
  assign or_981__in0[15:0] = in_1962[15:0];
  assign or_981__in1[15:0] = in_1963[15:0];
  assign reg_981__in[15:0] = or_981__out[15:0];
  assign or_983__in0[15:0] = in_1966[15:0];
  assign or_983__in1[15:0] = in_1967[15:0];
  assign reg_983__in[15:0] = or_983__out[15:0];
  assign or_985__in0[15:0] = in_1970[15:0];
  assign or_985__in1[15:0] = in_1971[15:0];
  assign reg_985__in[15:0] = or_985__out[15:0];
  assign or_987__in0[15:0] = in_1974[15:0];
  assign or_987__in1[15:0] = in_1975[15:0];
  assign reg_987__in[15:0] = or_987__out[15:0];
  assign or_989__in0[15:0] = in_1978[15:0];
  assign or_989__in1[15:0] = in_1979[15:0];
  assign reg_989__in[15:0] = or_989__out[15:0];
  assign or_99__in0[15:0] = in_198[15:0];
  assign or_99__in1[15:0] = in_199[15:0];
  assign reg_99__in[15:0] = or_99__out[15:0];
  assign or_991__in0[15:0] = in_1982[15:0];
  assign or_991__in1[15:0] = in_1983[15:0];
  assign reg_991__in[15:0] = or_991__out[15:0];
  assign or_993__in0[15:0] = in_1986[15:0];
  assign or_993__in1[15:0] = in_1987[15:0];
  assign reg_993__in[15:0] = or_993__out[15:0];
  assign or_995__in0[15:0] = in_1990[15:0];
  assign or_995__in1[15:0] = in_1991[15:0];
  assign reg_995__in[15:0] = or_995__out[15:0];
  assign or_997__in0[15:0] = in_1994[15:0];
  assign or_997__in1[15:0] = in_1995[15:0];
  assign reg_997__in[15:0] = or_997__out[15:0];
  assign or_999__in0[15:0] = in_1998[15:0];
  assign or_999__in1[15:0] = in_1999[15:0];
  assign reg_999__in[15:0] = or_999__out[15:0];
  assign reg_0__clk = clk;
  assign out_0[15:0] = reg_0__out[15:0];
  assign reg_1__clk = clk;
  assign out_1[15:0] = reg_1__out[15:0];
  assign reg_10__clk = clk;
  assign out_10[15:0] = reg_10__out[15:0];
  assign reg_100__clk = clk;
  assign out_100[15:0] = reg_100__out[15:0];
  assign reg_101__clk = clk;
  assign out_101[15:0] = reg_101__out[15:0];
  assign reg_102__clk = clk;
  assign out_102[15:0] = reg_102__out[15:0];
  assign reg_103__clk = clk;
  assign out_103[15:0] = reg_103__out[15:0];
  assign reg_104__clk = clk;
  assign out_104[15:0] = reg_104__out[15:0];
  assign reg_105__clk = clk;
  assign out_105[15:0] = reg_105__out[15:0];
  assign reg_106__clk = clk;
  assign out_106[15:0] = reg_106__out[15:0];
  assign reg_107__clk = clk;
  assign out_107[15:0] = reg_107__out[15:0];
  assign reg_108__clk = clk;
  assign out_108[15:0] = reg_108__out[15:0];
  assign reg_109__clk = clk;
  assign out_109[15:0] = reg_109__out[15:0];
  assign reg_11__clk = clk;
  assign out_11[15:0] = reg_11__out[15:0];
  assign reg_110__clk = clk;
  assign out_110[15:0] = reg_110__out[15:0];
  assign reg_111__clk = clk;
  assign out_111[15:0] = reg_111__out[15:0];
  assign reg_112__clk = clk;
  assign out_112[15:0] = reg_112__out[15:0];
  assign reg_113__clk = clk;
  assign out_113[15:0] = reg_113__out[15:0];
  assign reg_114__clk = clk;
  assign out_114[15:0] = reg_114__out[15:0];
  assign reg_115__clk = clk;
  assign out_115[15:0] = reg_115__out[15:0];
  assign reg_116__clk = clk;
  assign out_116[15:0] = reg_116__out[15:0];
  assign reg_117__clk = clk;
  assign out_117[15:0] = reg_117__out[15:0];
  assign reg_118__clk = clk;
  assign out_118[15:0] = reg_118__out[15:0];
  assign reg_119__clk = clk;
  assign out_119[15:0] = reg_119__out[15:0];
  assign reg_12__clk = clk;
  assign out_12[15:0] = reg_12__out[15:0];
  assign reg_120__clk = clk;
  assign out_120[15:0] = reg_120__out[15:0];
  assign reg_121__clk = clk;
  assign out_121[15:0] = reg_121__out[15:0];
  assign reg_122__clk = clk;
  assign out_122[15:0] = reg_122__out[15:0];
  assign reg_123__clk = clk;
  assign out_123[15:0] = reg_123__out[15:0];
  assign reg_124__clk = clk;
  assign out_124[15:0] = reg_124__out[15:0];
  assign reg_125__clk = clk;
  assign out_125[15:0] = reg_125__out[15:0];
  assign reg_126__clk = clk;
  assign out_126[15:0] = reg_126__out[15:0];
  assign reg_127__clk = clk;
  assign out_127[15:0] = reg_127__out[15:0];
  assign reg_128__clk = clk;
  assign out_128[15:0] = reg_128__out[15:0];
  assign reg_129__clk = clk;
  assign out_129[15:0] = reg_129__out[15:0];
  assign reg_13__clk = clk;
  assign out_13[15:0] = reg_13__out[15:0];
  assign reg_130__clk = clk;
  assign out_130[15:0] = reg_130__out[15:0];
  assign reg_131__clk = clk;
  assign out_131[15:0] = reg_131__out[15:0];
  assign reg_132__clk = clk;
  assign out_132[15:0] = reg_132__out[15:0];
  assign reg_133__clk = clk;
  assign out_133[15:0] = reg_133__out[15:0];
  assign reg_134__clk = clk;
  assign out_134[15:0] = reg_134__out[15:0];
  assign reg_135__clk = clk;
  assign out_135[15:0] = reg_135__out[15:0];
  assign reg_136__clk = clk;
  assign out_136[15:0] = reg_136__out[15:0];
  assign reg_137__clk = clk;
  assign out_137[15:0] = reg_137__out[15:0];
  assign reg_138__clk = clk;
  assign out_138[15:0] = reg_138__out[15:0];
  assign reg_139__clk = clk;
  assign out_139[15:0] = reg_139__out[15:0];
  assign reg_14__clk = clk;
  assign out_14[15:0] = reg_14__out[15:0];
  assign reg_140__clk = clk;
  assign out_140[15:0] = reg_140__out[15:0];
  assign reg_141__clk = clk;
  assign out_141[15:0] = reg_141__out[15:0];
  assign reg_142__clk = clk;
  assign out_142[15:0] = reg_142__out[15:0];
  assign reg_143__clk = clk;
  assign out_143[15:0] = reg_143__out[15:0];
  assign reg_144__clk = clk;
  assign out_144[15:0] = reg_144__out[15:0];
  assign reg_145__clk = clk;
  assign out_145[15:0] = reg_145__out[15:0];
  assign reg_146__clk = clk;
  assign out_146[15:0] = reg_146__out[15:0];
  assign reg_147__clk = clk;
  assign out_147[15:0] = reg_147__out[15:0];
  assign reg_148__clk = clk;
  assign out_148[15:0] = reg_148__out[15:0];
  assign reg_149__clk = clk;
  assign out_149[15:0] = reg_149__out[15:0];
  assign reg_15__clk = clk;
  assign out_15[15:0] = reg_15__out[15:0];
  assign reg_150__clk = clk;
  assign out_150[15:0] = reg_150__out[15:0];
  assign reg_151__clk = clk;
  assign out_151[15:0] = reg_151__out[15:0];
  assign reg_152__clk = clk;
  assign out_152[15:0] = reg_152__out[15:0];
  assign reg_153__clk = clk;
  assign out_153[15:0] = reg_153__out[15:0];
  assign reg_154__clk = clk;
  assign out_154[15:0] = reg_154__out[15:0];
  assign reg_155__clk = clk;
  assign out_155[15:0] = reg_155__out[15:0];
  assign reg_156__clk = clk;
  assign out_156[15:0] = reg_156__out[15:0];
  assign reg_157__clk = clk;
  assign out_157[15:0] = reg_157__out[15:0];
  assign reg_158__clk = clk;
  assign out_158[15:0] = reg_158__out[15:0];
  assign reg_159__clk = clk;
  assign out_159[15:0] = reg_159__out[15:0];
  assign reg_16__clk = clk;
  assign out_16[15:0] = reg_16__out[15:0];
  assign reg_160__clk = clk;
  assign out_160[15:0] = reg_160__out[15:0];
  assign reg_161__clk = clk;
  assign out_161[15:0] = reg_161__out[15:0];
  assign reg_162__clk = clk;
  assign out_162[15:0] = reg_162__out[15:0];
  assign reg_163__clk = clk;
  assign out_163[15:0] = reg_163__out[15:0];
  assign reg_164__clk = clk;
  assign out_164[15:0] = reg_164__out[15:0];
  assign reg_165__clk = clk;
  assign out_165[15:0] = reg_165__out[15:0];
  assign reg_166__clk = clk;
  assign out_166[15:0] = reg_166__out[15:0];
  assign reg_167__clk = clk;
  assign out_167[15:0] = reg_167__out[15:0];
  assign reg_168__clk = clk;
  assign out_168[15:0] = reg_168__out[15:0];
  assign reg_169__clk = clk;
  assign out_169[15:0] = reg_169__out[15:0];
  assign reg_17__clk = clk;
  assign out_17[15:0] = reg_17__out[15:0];
  assign reg_170__clk = clk;
  assign out_170[15:0] = reg_170__out[15:0];
  assign reg_171__clk = clk;
  assign out_171[15:0] = reg_171__out[15:0];
  assign reg_172__clk = clk;
  assign out_172[15:0] = reg_172__out[15:0];
  assign reg_173__clk = clk;
  assign out_173[15:0] = reg_173__out[15:0];
  assign reg_174__clk = clk;
  assign out_174[15:0] = reg_174__out[15:0];
  assign reg_175__clk = clk;
  assign out_175[15:0] = reg_175__out[15:0];
  assign reg_176__clk = clk;
  assign out_176[15:0] = reg_176__out[15:0];
  assign reg_177__clk = clk;
  assign out_177[15:0] = reg_177__out[15:0];
  assign reg_178__clk = clk;
  assign out_178[15:0] = reg_178__out[15:0];
  assign reg_179__clk = clk;
  assign out_179[15:0] = reg_179__out[15:0];
  assign reg_18__clk = clk;
  assign out_18[15:0] = reg_18__out[15:0];
  assign reg_180__clk = clk;
  assign out_180[15:0] = reg_180__out[15:0];
  assign reg_181__clk = clk;
  assign out_181[15:0] = reg_181__out[15:0];
  assign reg_182__clk = clk;
  assign out_182[15:0] = reg_182__out[15:0];
  assign reg_183__clk = clk;
  assign out_183[15:0] = reg_183__out[15:0];
  assign reg_184__clk = clk;
  assign out_184[15:0] = reg_184__out[15:0];
  assign reg_185__clk = clk;
  assign out_185[15:0] = reg_185__out[15:0];
  assign reg_186__clk = clk;
  assign out_186[15:0] = reg_186__out[15:0];
  assign reg_187__clk = clk;
  assign out_187[15:0] = reg_187__out[15:0];
  assign reg_188__clk = clk;
  assign out_188[15:0] = reg_188__out[15:0];
  assign reg_189__clk = clk;
  assign out_189[15:0] = reg_189__out[15:0];
  assign reg_19__clk = clk;
  assign out_19[15:0] = reg_19__out[15:0];
  assign reg_190__clk = clk;
  assign out_190[15:0] = reg_190__out[15:0];
  assign reg_191__clk = clk;
  assign out_191[15:0] = reg_191__out[15:0];
  assign reg_192__clk = clk;
  assign out_192[15:0] = reg_192__out[15:0];
  assign reg_193__clk = clk;
  assign out_193[15:0] = reg_193__out[15:0];
  assign reg_194__clk = clk;
  assign out_194[15:0] = reg_194__out[15:0];
  assign reg_195__clk = clk;
  assign out_195[15:0] = reg_195__out[15:0];
  assign reg_196__clk = clk;
  assign out_196[15:0] = reg_196__out[15:0];
  assign reg_197__clk = clk;
  assign out_197[15:0] = reg_197__out[15:0];
  assign reg_198__clk = clk;
  assign out_198[15:0] = reg_198__out[15:0];
  assign reg_199__clk = clk;
  assign out_199[15:0] = reg_199__out[15:0];
  assign reg_2__clk = clk;
  assign out_2[15:0] = reg_2__out[15:0];
  assign reg_20__clk = clk;
  assign out_20[15:0] = reg_20__out[15:0];
  assign reg_200__clk = clk;
  assign out_200[15:0] = reg_200__out[15:0];
  assign reg_201__clk = clk;
  assign out_201[15:0] = reg_201__out[15:0];
  assign reg_202__clk = clk;
  assign out_202[15:0] = reg_202__out[15:0];
  assign reg_203__clk = clk;
  assign out_203[15:0] = reg_203__out[15:0];
  assign reg_204__clk = clk;
  assign out_204[15:0] = reg_204__out[15:0];
  assign reg_205__clk = clk;
  assign out_205[15:0] = reg_205__out[15:0];
  assign reg_206__clk = clk;
  assign out_206[15:0] = reg_206__out[15:0];
  assign reg_207__clk = clk;
  assign out_207[15:0] = reg_207__out[15:0];
  assign reg_208__clk = clk;
  assign out_208[15:0] = reg_208__out[15:0];
  assign reg_209__clk = clk;
  assign out_209[15:0] = reg_209__out[15:0];
  assign reg_21__clk = clk;
  assign out_21[15:0] = reg_21__out[15:0];
  assign reg_210__clk = clk;
  assign out_210[15:0] = reg_210__out[15:0];
  assign reg_211__clk = clk;
  assign out_211[15:0] = reg_211__out[15:0];
  assign reg_212__clk = clk;
  assign out_212[15:0] = reg_212__out[15:0];
  assign reg_213__clk = clk;
  assign out_213[15:0] = reg_213__out[15:0];
  assign reg_214__clk = clk;
  assign out_214[15:0] = reg_214__out[15:0];
  assign reg_215__clk = clk;
  assign out_215[15:0] = reg_215__out[15:0];
  assign reg_216__clk = clk;
  assign out_216[15:0] = reg_216__out[15:0];
  assign reg_217__clk = clk;
  assign out_217[15:0] = reg_217__out[15:0];
  assign reg_218__clk = clk;
  assign out_218[15:0] = reg_218__out[15:0];
  assign reg_219__clk = clk;
  assign out_219[15:0] = reg_219__out[15:0];
  assign reg_22__clk = clk;
  assign out_22[15:0] = reg_22__out[15:0];
  assign reg_220__clk = clk;
  assign out_220[15:0] = reg_220__out[15:0];
  assign reg_221__clk = clk;
  assign out_221[15:0] = reg_221__out[15:0];
  assign reg_222__clk = clk;
  assign out_222[15:0] = reg_222__out[15:0];
  assign reg_223__clk = clk;
  assign out_223[15:0] = reg_223__out[15:0];
  assign reg_224__clk = clk;
  assign out_224[15:0] = reg_224__out[15:0];
  assign reg_225__clk = clk;
  assign out_225[15:0] = reg_225__out[15:0];
  assign reg_226__clk = clk;
  assign out_226[15:0] = reg_226__out[15:0];
  assign reg_227__clk = clk;
  assign out_227[15:0] = reg_227__out[15:0];
  assign reg_228__clk = clk;
  assign out_228[15:0] = reg_228__out[15:0];
  assign reg_229__clk = clk;
  assign out_229[15:0] = reg_229__out[15:0];
  assign reg_23__clk = clk;
  assign out_23[15:0] = reg_23__out[15:0];
  assign reg_230__clk = clk;
  assign out_230[15:0] = reg_230__out[15:0];
  assign reg_231__clk = clk;
  assign out_231[15:0] = reg_231__out[15:0];
  assign reg_232__clk = clk;
  assign out_232[15:0] = reg_232__out[15:0];
  assign reg_233__clk = clk;
  assign out_233[15:0] = reg_233__out[15:0];
  assign reg_234__clk = clk;
  assign out_234[15:0] = reg_234__out[15:0];
  assign reg_235__clk = clk;
  assign out_235[15:0] = reg_235__out[15:0];
  assign reg_236__clk = clk;
  assign out_236[15:0] = reg_236__out[15:0];
  assign reg_237__clk = clk;
  assign out_237[15:0] = reg_237__out[15:0];
  assign reg_238__clk = clk;
  assign out_238[15:0] = reg_238__out[15:0];
  assign reg_239__clk = clk;
  assign out_239[15:0] = reg_239__out[15:0];
  assign reg_24__clk = clk;
  assign out_24[15:0] = reg_24__out[15:0];
  assign reg_240__clk = clk;
  assign out_240[15:0] = reg_240__out[15:0];
  assign reg_241__clk = clk;
  assign out_241[15:0] = reg_241__out[15:0];
  assign reg_242__clk = clk;
  assign out_242[15:0] = reg_242__out[15:0];
  assign reg_243__clk = clk;
  assign out_243[15:0] = reg_243__out[15:0];
  assign reg_244__clk = clk;
  assign out_244[15:0] = reg_244__out[15:0];
  assign reg_245__clk = clk;
  assign out_245[15:0] = reg_245__out[15:0];
  assign reg_246__clk = clk;
  assign out_246[15:0] = reg_246__out[15:0];
  assign reg_247__clk = clk;
  assign out_247[15:0] = reg_247__out[15:0];
  assign reg_248__clk = clk;
  assign out_248[15:0] = reg_248__out[15:0];
  assign reg_249__clk = clk;
  assign out_249[15:0] = reg_249__out[15:0];
  assign reg_25__clk = clk;
  assign out_25[15:0] = reg_25__out[15:0];
  assign reg_250__clk = clk;
  assign out_250[15:0] = reg_250__out[15:0];
  assign reg_251__clk = clk;
  assign out_251[15:0] = reg_251__out[15:0];
  assign reg_252__clk = clk;
  assign out_252[15:0] = reg_252__out[15:0];
  assign reg_253__clk = clk;
  assign out_253[15:0] = reg_253__out[15:0];
  assign reg_254__clk = clk;
  assign out_254[15:0] = reg_254__out[15:0];
  assign reg_255__clk = clk;
  assign out_255[15:0] = reg_255__out[15:0];
  assign reg_256__clk = clk;
  assign out_256[15:0] = reg_256__out[15:0];
  assign reg_257__clk = clk;
  assign out_257[15:0] = reg_257__out[15:0];
  assign reg_258__clk = clk;
  assign out_258[15:0] = reg_258__out[15:0];
  assign reg_259__clk = clk;
  assign out_259[15:0] = reg_259__out[15:0];
  assign reg_26__clk = clk;
  assign out_26[15:0] = reg_26__out[15:0];
  assign reg_260__clk = clk;
  assign out_260[15:0] = reg_260__out[15:0];
  assign reg_261__clk = clk;
  assign out_261[15:0] = reg_261__out[15:0];
  assign reg_262__clk = clk;
  assign out_262[15:0] = reg_262__out[15:0];
  assign reg_263__clk = clk;
  assign out_263[15:0] = reg_263__out[15:0];
  assign reg_264__clk = clk;
  assign out_264[15:0] = reg_264__out[15:0];
  assign reg_265__clk = clk;
  assign out_265[15:0] = reg_265__out[15:0];
  assign reg_266__clk = clk;
  assign out_266[15:0] = reg_266__out[15:0];
  assign reg_267__clk = clk;
  assign out_267[15:0] = reg_267__out[15:0];
  assign reg_268__clk = clk;
  assign out_268[15:0] = reg_268__out[15:0];
  assign reg_269__clk = clk;
  assign out_269[15:0] = reg_269__out[15:0];
  assign reg_27__clk = clk;
  assign out_27[15:0] = reg_27__out[15:0];
  assign reg_270__clk = clk;
  assign out_270[15:0] = reg_270__out[15:0];
  assign reg_271__clk = clk;
  assign out_271[15:0] = reg_271__out[15:0];
  assign reg_272__clk = clk;
  assign out_272[15:0] = reg_272__out[15:0];
  assign reg_273__clk = clk;
  assign out_273[15:0] = reg_273__out[15:0];
  assign reg_274__clk = clk;
  assign out_274[15:0] = reg_274__out[15:0];
  assign reg_275__clk = clk;
  assign out_275[15:0] = reg_275__out[15:0];
  assign reg_276__clk = clk;
  assign out_276[15:0] = reg_276__out[15:0];
  assign reg_277__clk = clk;
  assign out_277[15:0] = reg_277__out[15:0];
  assign reg_278__clk = clk;
  assign out_278[15:0] = reg_278__out[15:0];
  assign reg_279__clk = clk;
  assign out_279[15:0] = reg_279__out[15:0];
  assign reg_28__clk = clk;
  assign out_28[15:0] = reg_28__out[15:0];
  assign reg_280__clk = clk;
  assign out_280[15:0] = reg_280__out[15:0];
  assign reg_281__clk = clk;
  assign out_281[15:0] = reg_281__out[15:0];
  assign reg_282__clk = clk;
  assign out_282[15:0] = reg_282__out[15:0];
  assign reg_283__clk = clk;
  assign out_283[15:0] = reg_283__out[15:0];
  assign reg_284__clk = clk;
  assign out_284[15:0] = reg_284__out[15:0];
  assign reg_285__clk = clk;
  assign out_285[15:0] = reg_285__out[15:0];
  assign reg_286__clk = clk;
  assign out_286[15:0] = reg_286__out[15:0];
  assign reg_287__clk = clk;
  assign out_287[15:0] = reg_287__out[15:0];
  assign reg_288__clk = clk;
  assign out_288[15:0] = reg_288__out[15:0];
  assign reg_289__clk = clk;
  assign out_289[15:0] = reg_289__out[15:0];
  assign reg_29__clk = clk;
  assign out_29[15:0] = reg_29__out[15:0];
  assign reg_290__clk = clk;
  assign out_290[15:0] = reg_290__out[15:0];
  assign reg_291__clk = clk;
  assign out_291[15:0] = reg_291__out[15:0];
  assign reg_292__clk = clk;
  assign out_292[15:0] = reg_292__out[15:0];
  assign reg_293__clk = clk;
  assign out_293[15:0] = reg_293__out[15:0];
  assign reg_294__clk = clk;
  assign out_294[15:0] = reg_294__out[15:0];
  assign reg_295__clk = clk;
  assign out_295[15:0] = reg_295__out[15:0];
  assign reg_296__clk = clk;
  assign out_296[15:0] = reg_296__out[15:0];
  assign reg_297__clk = clk;
  assign out_297[15:0] = reg_297__out[15:0];
  assign reg_298__clk = clk;
  assign out_298[15:0] = reg_298__out[15:0];
  assign reg_299__clk = clk;
  assign out_299[15:0] = reg_299__out[15:0];
  assign reg_3__clk = clk;
  assign out_3[15:0] = reg_3__out[15:0];
  assign reg_30__clk = clk;
  assign out_30[15:0] = reg_30__out[15:0];
  assign reg_300__clk = clk;
  assign out_300[15:0] = reg_300__out[15:0];
  assign reg_301__clk = clk;
  assign out_301[15:0] = reg_301__out[15:0];
  assign reg_302__clk = clk;
  assign out_302[15:0] = reg_302__out[15:0];
  assign reg_303__clk = clk;
  assign out_303[15:0] = reg_303__out[15:0];
  assign reg_304__clk = clk;
  assign out_304[15:0] = reg_304__out[15:0];
  assign reg_305__clk = clk;
  assign out_305[15:0] = reg_305__out[15:0];
  assign reg_306__clk = clk;
  assign out_306[15:0] = reg_306__out[15:0];
  assign reg_307__clk = clk;
  assign out_307[15:0] = reg_307__out[15:0];
  assign reg_308__clk = clk;
  assign out_308[15:0] = reg_308__out[15:0];
  assign reg_309__clk = clk;
  assign out_309[15:0] = reg_309__out[15:0];
  assign reg_31__clk = clk;
  assign out_31[15:0] = reg_31__out[15:0];
  assign reg_310__clk = clk;
  assign out_310[15:0] = reg_310__out[15:0];
  assign reg_311__clk = clk;
  assign out_311[15:0] = reg_311__out[15:0];
  assign reg_312__clk = clk;
  assign out_312[15:0] = reg_312__out[15:0];
  assign reg_313__clk = clk;
  assign out_313[15:0] = reg_313__out[15:0];
  assign reg_314__clk = clk;
  assign out_314[15:0] = reg_314__out[15:0];
  assign reg_315__clk = clk;
  assign out_315[15:0] = reg_315__out[15:0];
  assign reg_316__clk = clk;
  assign out_316[15:0] = reg_316__out[15:0];
  assign reg_317__clk = clk;
  assign out_317[15:0] = reg_317__out[15:0];
  assign reg_318__clk = clk;
  assign out_318[15:0] = reg_318__out[15:0];
  assign reg_319__clk = clk;
  assign out_319[15:0] = reg_319__out[15:0];
  assign reg_32__clk = clk;
  assign out_32[15:0] = reg_32__out[15:0];
  assign reg_320__clk = clk;
  assign out_320[15:0] = reg_320__out[15:0];
  assign reg_321__clk = clk;
  assign out_321[15:0] = reg_321__out[15:0];
  assign reg_322__clk = clk;
  assign out_322[15:0] = reg_322__out[15:0];
  assign reg_323__clk = clk;
  assign out_323[15:0] = reg_323__out[15:0];
  assign reg_324__clk = clk;
  assign out_324[15:0] = reg_324__out[15:0];
  assign reg_325__clk = clk;
  assign out_325[15:0] = reg_325__out[15:0];
  assign reg_326__clk = clk;
  assign out_326[15:0] = reg_326__out[15:0];
  assign reg_327__clk = clk;
  assign out_327[15:0] = reg_327__out[15:0];
  assign reg_328__clk = clk;
  assign out_328[15:0] = reg_328__out[15:0];
  assign reg_329__clk = clk;
  assign out_329[15:0] = reg_329__out[15:0];
  assign reg_33__clk = clk;
  assign out_33[15:0] = reg_33__out[15:0];
  assign reg_330__clk = clk;
  assign out_330[15:0] = reg_330__out[15:0];
  assign reg_331__clk = clk;
  assign out_331[15:0] = reg_331__out[15:0];
  assign reg_332__clk = clk;
  assign out_332[15:0] = reg_332__out[15:0];
  assign reg_333__clk = clk;
  assign out_333[15:0] = reg_333__out[15:0];
  assign reg_334__clk = clk;
  assign out_334[15:0] = reg_334__out[15:0];
  assign reg_335__clk = clk;
  assign out_335[15:0] = reg_335__out[15:0];
  assign reg_336__clk = clk;
  assign out_336[15:0] = reg_336__out[15:0];
  assign reg_337__clk = clk;
  assign out_337[15:0] = reg_337__out[15:0];
  assign reg_338__clk = clk;
  assign out_338[15:0] = reg_338__out[15:0];
  assign reg_339__clk = clk;
  assign out_339[15:0] = reg_339__out[15:0];
  assign reg_34__clk = clk;
  assign out_34[15:0] = reg_34__out[15:0];
  assign reg_340__clk = clk;
  assign out_340[15:0] = reg_340__out[15:0];
  assign reg_341__clk = clk;
  assign out_341[15:0] = reg_341__out[15:0];
  assign reg_342__clk = clk;
  assign out_342[15:0] = reg_342__out[15:0];
  assign reg_343__clk = clk;
  assign out_343[15:0] = reg_343__out[15:0];
  assign reg_344__clk = clk;
  assign out_344[15:0] = reg_344__out[15:0];
  assign reg_345__clk = clk;
  assign out_345[15:0] = reg_345__out[15:0];
  assign reg_346__clk = clk;
  assign out_346[15:0] = reg_346__out[15:0];
  assign reg_347__clk = clk;
  assign out_347[15:0] = reg_347__out[15:0];
  assign reg_348__clk = clk;
  assign out_348[15:0] = reg_348__out[15:0];
  assign reg_349__clk = clk;
  assign out_349[15:0] = reg_349__out[15:0];
  assign reg_35__clk = clk;
  assign out_35[15:0] = reg_35__out[15:0];
  assign reg_350__clk = clk;
  assign out_350[15:0] = reg_350__out[15:0];
  assign reg_351__clk = clk;
  assign out_351[15:0] = reg_351__out[15:0];
  assign reg_352__clk = clk;
  assign out_352[15:0] = reg_352__out[15:0];
  assign reg_353__clk = clk;
  assign out_353[15:0] = reg_353__out[15:0];
  assign reg_354__clk = clk;
  assign out_354[15:0] = reg_354__out[15:0];
  assign reg_355__clk = clk;
  assign out_355[15:0] = reg_355__out[15:0];
  assign reg_356__clk = clk;
  assign out_356[15:0] = reg_356__out[15:0];
  assign reg_357__clk = clk;
  assign out_357[15:0] = reg_357__out[15:0];
  assign reg_358__clk = clk;
  assign out_358[15:0] = reg_358__out[15:0];
  assign reg_359__clk = clk;
  assign out_359[15:0] = reg_359__out[15:0];
  assign reg_36__clk = clk;
  assign out_36[15:0] = reg_36__out[15:0];
  assign reg_360__clk = clk;
  assign out_360[15:0] = reg_360__out[15:0];
  assign reg_361__clk = clk;
  assign out_361[15:0] = reg_361__out[15:0];
  assign reg_362__clk = clk;
  assign out_362[15:0] = reg_362__out[15:0];
  assign reg_363__clk = clk;
  assign out_363[15:0] = reg_363__out[15:0];
  assign reg_364__clk = clk;
  assign out_364[15:0] = reg_364__out[15:0];
  assign reg_365__clk = clk;
  assign out_365[15:0] = reg_365__out[15:0];
  assign reg_366__clk = clk;
  assign out_366[15:0] = reg_366__out[15:0];
  assign reg_367__clk = clk;
  assign out_367[15:0] = reg_367__out[15:0];
  assign reg_368__clk = clk;
  assign out_368[15:0] = reg_368__out[15:0];
  assign reg_369__clk = clk;
  assign out_369[15:0] = reg_369__out[15:0];
  assign reg_37__clk = clk;
  assign out_37[15:0] = reg_37__out[15:0];
  assign reg_370__clk = clk;
  assign out_370[15:0] = reg_370__out[15:0];
  assign reg_371__clk = clk;
  assign out_371[15:0] = reg_371__out[15:0];
  assign reg_372__clk = clk;
  assign out_372[15:0] = reg_372__out[15:0];
  assign reg_373__clk = clk;
  assign out_373[15:0] = reg_373__out[15:0];
  assign reg_374__clk = clk;
  assign out_374[15:0] = reg_374__out[15:0];
  assign reg_375__clk = clk;
  assign out_375[15:0] = reg_375__out[15:0];
  assign reg_376__clk = clk;
  assign out_376[15:0] = reg_376__out[15:0];
  assign reg_377__clk = clk;
  assign out_377[15:0] = reg_377__out[15:0];
  assign reg_378__clk = clk;
  assign out_378[15:0] = reg_378__out[15:0];
  assign reg_379__clk = clk;
  assign out_379[15:0] = reg_379__out[15:0];
  assign reg_38__clk = clk;
  assign out_38[15:0] = reg_38__out[15:0];
  assign reg_380__clk = clk;
  assign out_380[15:0] = reg_380__out[15:0];
  assign reg_381__clk = clk;
  assign out_381[15:0] = reg_381__out[15:0];
  assign reg_382__clk = clk;
  assign out_382[15:0] = reg_382__out[15:0];
  assign reg_383__clk = clk;
  assign out_383[15:0] = reg_383__out[15:0];
  assign reg_384__clk = clk;
  assign out_384[15:0] = reg_384__out[15:0];
  assign reg_385__clk = clk;
  assign out_385[15:0] = reg_385__out[15:0];
  assign reg_386__clk = clk;
  assign out_386[15:0] = reg_386__out[15:0];
  assign reg_387__clk = clk;
  assign out_387[15:0] = reg_387__out[15:0];
  assign reg_388__clk = clk;
  assign out_388[15:0] = reg_388__out[15:0];
  assign reg_389__clk = clk;
  assign out_389[15:0] = reg_389__out[15:0];
  assign reg_39__clk = clk;
  assign out_39[15:0] = reg_39__out[15:0];
  assign reg_390__clk = clk;
  assign out_390[15:0] = reg_390__out[15:0];
  assign reg_391__clk = clk;
  assign out_391[15:0] = reg_391__out[15:0];
  assign reg_392__clk = clk;
  assign out_392[15:0] = reg_392__out[15:0];
  assign reg_393__clk = clk;
  assign out_393[15:0] = reg_393__out[15:0];
  assign reg_394__clk = clk;
  assign out_394[15:0] = reg_394__out[15:0];
  assign reg_395__clk = clk;
  assign out_395[15:0] = reg_395__out[15:0];
  assign reg_396__clk = clk;
  assign out_396[15:0] = reg_396__out[15:0];
  assign reg_397__clk = clk;
  assign out_397[15:0] = reg_397__out[15:0];
  assign reg_398__clk = clk;
  assign out_398[15:0] = reg_398__out[15:0];
  assign reg_399__clk = clk;
  assign out_399[15:0] = reg_399__out[15:0];
  assign reg_4__clk = clk;
  assign out_4[15:0] = reg_4__out[15:0];
  assign reg_40__clk = clk;
  assign out_40[15:0] = reg_40__out[15:0];
  assign reg_400__clk = clk;
  assign out_400[15:0] = reg_400__out[15:0];
  assign reg_401__clk = clk;
  assign out_401[15:0] = reg_401__out[15:0];
  assign reg_402__clk = clk;
  assign out_402[15:0] = reg_402__out[15:0];
  assign reg_403__clk = clk;
  assign out_403[15:0] = reg_403__out[15:0];
  assign reg_404__clk = clk;
  assign out_404[15:0] = reg_404__out[15:0];
  assign reg_405__clk = clk;
  assign out_405[15:0] = reg_405__out[15:0];
  assign reg_406__clk = clk;
  assign out_406[15:0] = reg_406__out[15:0];
  assign reg_407__clk = clk;
  assign out_407[15:0] = reg_407__out[15:0];
  assign reg_408__clk = clk;
  assign out_408[15:0] = reg_408__out[15:0];
  assign reg_409__clk = clk;
  assign out_409[15:0] = reg_409__out[15:0];
  assign reg_41__clk = clk;
  assign out_41[15:0] = reg_41__out[15:0];
  assign reg_410__clk = clk;
  assign out_410[15:0] = reg_410__out[15:0];
  assign reg_411__clk = clk;
  assign out_411[15:0] = reg_411__out[15:0];
  assign reg_412__clk = clk;
  assign out_412[15:0] = reg_412__out[15:0];
  assign reg_413__clk = clk;
  assign out_413[15:0] = reg_413__out[15:0];
  assign reg_414__clk = clk;
  assign out_414[15:0] = reg_414__out[15:0];
  assign reg_415__clk = clk;
  assign out_415[15:0] = reg_415__out[15:0];
  assign reg_416__clk = clk;
  assign out_416[15:0] = reg_416__out[15:0];
  assign reg_417__clk = clk;
  assign out_417[15:0] = reg_417__out[15:0];
  assign reg_418__clk = clk;
  assign out_418[15:0] = reg_418__out[15:0];
  assign reg_419__clk = clk;
  assign out_419[15:0] = reg_419__out[15:0];
  assign reg_42__clk = clk;
  assign out_42[15:0] = reg_42__out[15:0];
  assign reg_420__clk = clk;
  assign out_420[15:0] = reg_420__out[15:0];
  assign reg_421__clk = clk;
  assign out_421[15:0] = reg_421__out[15:0];
  assign reg_422__clk = clk;
  assign out_422[15:0] = reg_422__out[15:0];
  assign reg_423__clk = clk;
  assign out_423[15:0] = reg_423__out[15:0];
  assign reg_424__clk = clk;
  assign out_424[15:0] = reg_424__out[15:0];
  assign reg_425__clk = clk;
  assign out_425[15:0] = reg_425__out[15:0];
  assign reg_426__clk = clk;
  assign out_426[15:0] = reg_426__out[15:0];
  assign reg_427__clk = clk;
  assign out_427[15:0] = reg_427__out[15:0];
  assign reg_428__clk = clk;
  assign out_428[15:0] = reg_428__out[15:0];
  assign reg_429__clk = clk;
  assign out_429[15:0] = reg_429__out[15:0];
  assign reg_43__clk = clk;
  assign out_43[15:0] = reg_43__out[15:0];
  assign reg_430__clk = clk;
  assign out_430[15:0] = reg_430__out[15:0];
  assign reg_431__clk = clk;
  assign out_431[15:0] = reg_431__out[15:0];
  assign reg_432__clk = clk;
  assign out_432[15:0] = reg_432__out[15:0];
  assign reg_433__clk = clk;
  assign out_433[15:0] = reg_433__out[15:0];
  assign reg_434__clk = clk;
  assign out_434[15:0] = reg_434__out[15:0];
  assign reg_435__clk = clk;
  assign out_435[15:0] = reg_435__out[15:0];
  assign reg_436__clk = clk;
  assign out_436[15:0] = reg_436__out[15:0];
  assign reg_437__clk = clk;
  assign out_437[15:0] = reg_437__out[15:0];
  assign reg_438__clk = clk;
  assign out_438[15:0] = reg_438__out[15:0];
  assign reg_439__clk = clk;
  assign out_439[15:0] = reg_439__out[15:0];
  assign reg_44__clk = clk;
  assign out_44[15:0] = reg_44__out[15:0];
  assign reg_440__clk = clk;
  assign out_440[15:0] = reg_440__out[15:0];
  assign reg_441__clk = clk;
  assign out_441[15:0] = reg_441__out[15:0];
  assign reg_442__clk = clk;
  assign out_442[15:0] = reg_442__out[15:0];
  assign reg_443__clk = clk;
  assign out_443[15:0] = reg_443__out[15:0];
  assign reg_444__clk = clk;
  assign out_444[15:0] = reg_444__out[15:0];
  assign reg_445__clk = clk;
  assign out_445[15:0] = reg_445__out[15:0];
  assign reg_446__clk = clk;
  assign out_446[15:0] = reg_446__out[15:0];
  assign reg_447__clk = clk;
  assign out_447[15:0] = reg_447__out[15:0];
  assign reg_448__clk = clk;
  assign out_448[15:0] = reg_448__out[15:0];
  assign reg_449__clk = clk;
  assign out_449[15:0] = reg_449__out[15:0];
  assign reg_45__clk = clk;
  assign out_45[15:0] = reg_45__out[15:0];
  assign reg_450__clk = clk;
  assign out_450[15:0] = reg_450__out[15:0];
  assign reg_451__clk = clk;
  assign out_451[15:0] = reg_451__out[15:0];
  assign reg_452__clk = clk;
  assign out_452[15:0] = reg_452__out[15:0];
  assign reg_453__clk = clk;
  assign out_453[15:0] = reg_453__out[15:0];
  assign reg_454__clk = clk;
  assign out_454[15:0] = reg_454__out[15:0];
  assign reg_455__clk = clk;
  assign out_455[15:0] = reg_455__out[15:0];
  assign reg_456__clk = clk;
  assign out_456[15:0] = reg_456__out[15:0];
  assign reg_457__clk = clk;
  assign out_457[15:0] = reg_457__out[15:0];
  assign reg_458__clk = clk;
  assign out_458[15:0] = reg_458__out[15:0];
  assign reg_459__clk = clk;
  assign out_459[15:0] = reg_459__out[15:0];
  assign reg_46__clk = clk;
  assign out_46[15:0] = reg_46__out[15:0];
  assign reg_460__clk = clk;
  assign out_460[15:0] = reg_460__out[15:0];
  assign reg_461__clk = clk;
  assign out_461[15:0] = reg_461__out[15:0];
  assign reg_462__clk = clk;
  assign out_462[15:0] = reg_462__out[15:0];
  assign reg_463__clk = clk;
  assign out_463[15:0] = reg_463__out[15:0];
  assign reg_464__clk = clk;
  assign out_464[15:0] = reg_464__out[15:0];
  assign reg_465__clk = clk;
  assign out_465[15:0] = reg_465__out[15:0];
  assign reg_466__clk = clk;
  assign out_466[15:0] = reg_466__out[15:0];
  assign reg_467__clk = clk;
  assign out_467[15:0] = reg_467__out[15:0];
  assign reg_468__clk = clk;
  assign out_468[15:0] = reg_468__out[15:0];
  assign reg_469__clk = clk;
  assign out_469[15:0] = reg_469__out[15:0];
  assign reg_47__clk = clk;
  assign out_47[15:0] = reg_47__out[15:0];
  assign reg_470__clk = clk;
  assign out_470[15:0] = reg_470__out[15:0];
  assign reg_471__clk = clk;
  assign out_471[15:0] = reg_471__out[15:0];
  assign reg_472__clk = clk;
  assign out_472[15:0] = reg_472__out[15:0];
  assign reg_473__clk = clk;
  assign out_473[15:0] = reg_473__out[15:0];
  assign reg_474__clk = clk;
  assign out_474[15:0] = reg_474__out[15:0];
  assign reg_475__clk = clk;
  assign out_475[15:0] = reg_475__out[15:0];
  assign reg_476__clk = clk;
  assign out_476[15:0] = reg_476__out[15:0];
  assign reg_477__clk = clk;
  assign out_477[15:0] = reg_477__out[15:0];
  assign reg_478__clk = clk;
  assign out_478[15:0] = reg_478__out[15:0];
  assign reg_479__clk = clk;
  assign out_479[15:0] = reg_479__out[15:0];
  assign reg_48__clk = clk;
  assign out_48[15:0] = reg_48__out[15:0];
  assign reg_480__clk = clk;
  assign out_480[15:0] = reg_480__out[15:0];
  assign reg_481__clk = clk;
  assign out_481[15:0] = reg_481__out[15:0];
  assign reg_482__clk = clk;
  assign out_482[15:0] = reg_482__out[15:0];
  assign reg_483__clk = clk;
  assign out_483[15:0] = reg_483__out[15:0];
  assign reg_484__clk = clk;
  assign out_484[15:0] = reg_484__out[15:0];
  assign reg_485__clk = clk;
  assign out_485[15:0] = reg_485__out[15:0];
  assign reg_486__clk = clk;
  assign out_486[15:0] = reg_486__out[15:0];
  assign reg_487__clk = clk;
  assign out_487[15:0] = reg_487__out[15:0];
  assign reg_488__clk = clk;
  assign out_488[15:0] = reg_488__out[15:0];
  assign reg_489__clk = clk;
  assign out_489[15:0] = reg_489__out[15:0];
  assign reg_49__clk = clk;
  assign out_49[15:0] = reg_49__out[15:0];
  assign reg_490__clk = clk;
  assign out_490[15:0] = reg_490__out[15:0];
  assign reg_491__clk = clk;
  assign out_491[15:0] = reg_491__out[15:0];
  assign reg_492__clk = clk;
  assign out_492[15:0] = reg_492__out[15:0];
  assign reg_493__clk = clk;
  assign out_493[15:0] = reg_493__out[15:0];
  assign reg_494__clk = clk;
  assign out_494[15:0] = reg_494__out[15:0];
  assign reg_495__clk = clk;
  assign out_495[15:0] = reg_495__out[15:0];
  assign reg_496__clk = clk;
  assign out_496[15:0] = reg_496__out[15:0];
  assign reg_497__clk = clk;
  assign out_497[15:0] = reg_497__out[15:0];
  assign reg_498__clk = clk;
  assign out_498[15:0] = reg_498__out[15:0];
  assign reg_499__clk = clk;
  assign out_499[15:0] = reg_499__out[15:0];
  assign reg_5__clk = clk;
  assign out_5[15:0] = reg_5__out[15:0];
  assign reg_50__clk = clk;
  assign out_50[15:0] = reg_50__out[15:0];
  assign reg_500__clk = clk;
  assign out_500[15:0] = reg_500__out[15:0];
  assign reg_501__clk = clk;
  assign out_501[15:0] = reg_501__out[15:0];
  assign reg_502__clk = clk;
  assign out_502[15:0] = reg_502__out[15:0];
  assign reg_503__clk = clk;
  assign out_503[15:0] = reg_503__out[15:0];
  assign reg_504__clk = clk;
  assign out_504[15:0] = reg_504__out[15:0];
  assign reg_505__clk = clk;
  assign out_505[15:0] = reg_505__out[15:0];
  assign reg_506__clk = clk;
  assign out_506[15:0] = reg_506__out[15:0];
  assign reg_507__clk = clk;
  assign out_507[15:0] = reg_507__out[15:0];
  assign reg_508__clk = clk;
  assign out_508[15:0] = reg_508__out[15:0];
  assign reg_509__clk = clk;
  assign out_509[15:0] = reg_509__out[15:0];
  assign reg_51__clk = clk;
  assign out_51[15:0] = reg_51__out[15:0];
  assign reg_510__clk = clk;
  assign out_510[15:0] = reg_510__out[15:0];
  assign reg_511__clk = clk;
  assign out_511[15:0] = reg_511__out[15:0];
  assign reg_512__clk = clk;
  assign out_512[15:0] = reg_512__out[15:0];
  assign reg_513__clk = clk;
  assign out_513[15:0] = reg_513__out[15:0];
  assign reg_514__clk = clk;
  assign out_514[15:0] = reg_514__out[15:0];
  assign reg_515__clk = clk;
  assign out_515[15:0] = reg_515__out[15:0];
  assign reg_516__clk = clk;
  assign out_516[15:0] = reg_516__out[15:0];
  assign reg_517__clk = clk;
  assign out_517[15:0] = reg_517__out[15:0];
  assign reg_518__clk = clk;
  assign out_518[15:0] = reg_518__out[15:0];
  assign reg_519__clk = clk;
  assign out_519[15:0] = reg_519__out[15:0];
  assign reg_52__clk = clk;
  assign out_52[15:0] = reg_52__out[15:0];
  assign reg_520__clk = clk;
  assign out_520[15:0] = reg_520__out[15:0];
  assign reg_521__clk = clk;
  assign out_521[15:0] = reg_521__out[15:0];
  assign reg_522__clk = clk;
  assign out_522[15:0] = reg_522__out[15:0];
  assign reg_523__clk = clk;
  assign out_523[15:0] = reg_523__out[15:0];
  assign reg_524__clk = clk;
  assign out_524[15:0] = reg_524__out[15:0];
  assign reg_525__clk = clk;
  assign out_525[15:0] = reg_525__out[15:0];
  assign reg_526__clk = clk;
  assign out_526[15:0] = reg_526__out[15:0];
  assign reg_527__clk = clk;
  assign out_527[15:0] = reg_527__out[15:0];
  assign reg_528__clk = clk;
  assign out_528[15:0] = reg_528__out[15:0];
  assign reg_529__clk = clk;
  assign out_529[15:0] = reg_529__out[15:0];
  assign reg_53__clk = clk;
  assign out_53[15:0] = reg_53__out[15:0];
  assign reg_530__clk = clk;
  assign out_530[15:0] = reg_530__out[15:0];
  assign reg_531__clk = clk;
  assign out_531[15:0] = reg_531__out[15:0];
  assign reg_532__clk = clk;
  assign out_532[15:0] = reg_532__out[15:0];
  assign reg_533__clk = clk;
  assign out_533[15:0] = reg_533__out[15:0];
  assign reg_534__clk = clk;
  assign out_534[15:0] = reg_534__out[15:0];
  assign reg_535__clk = clk;
  assign out_535[15:0] = reg_535__out[15:0];
  assign reg_536__clk = clk;
  assign out_536[15:0] = reg_536__out[15:0];
  assign reg_537__clk = clk;
  assign out_537[15:0] = reg_537__out[15:0];
  assign reg_538__clk = clk;
  assign out_538[15:0] = reg_538__out[15:0];
  assign reg_539__clk = clk;
  assign out_539[15:0] = reg_539__out[15:0];
  assign reg_54__clk = clk;
  assign out_54[15:0] = reg_54__out[15:0];
  assign reg_540__clk = clk;
  assign out_540[15:0] = reg_540__out[15:0];
  assign reg_541__clk = clk;
  assign out_541[15:0] = reg_541__out[15:0];
  assign reg_542__clk = clk;
  assign out_542[15:0] = reg_542__out[15:0];
  assign reg_543__clk = clk;
  assign out_543[15:0] = reg_543__out[15:0];
  assign reg_544__clk = clk;
  assign out_544[15:0] = reg_544__out[15:0];
  assign reg_545__clk = clk;
  assign out_545[15:0] = reg_545__out[15:0];
  assign reg_546__clk = clk;
  assign out_546[15:0] = reg_546__out[15:0];
  assign reg_547__clk = clk;
  assign out_547[15:0] = reg_547__out[15:0];
  assign reg_548__clk = clk;
  assign out_548[15:0] = reg_548__out[15:0];
  assign reg_549__clk = clk;
  assign out_549[15:0] = reg_549__out[15:0];
  assign reg_55__clk = clk;
  assign out_55[15:0] = reg_55__out[15:0];
  assign reg_550__clk = clk;
  assign out_550[15:0] = reg_550__out[15:0];
  assign reg_551__clk = clk;
  assign out_551[15:0] = reg_551__out[15:0];
  assign reg_552__clk = clk;
  assign out_552[15:0] = reg_552__out[15:0];
  assign reg_553__clk = clk;
  assign out_553[15:0] = reg_553__out[15:0];
  assign reg_554__clk = clk;
  assign out_554[15:0] = reg_554__out[15:0];
  assign reg_555__clk = clk;
  assign out_555[15:0] = reg_555__out[15:0];
  assign reg_556__clk = clk;
  assign out_556[15:0] = reg_556__out[15:0];
  assign reg_557__clk = clk;
  assign out_557[15:0] = reg_557__out[15:0];
  assign reg_558__clk = clk;
  assign out_558[15:0] = reg_558__out[15:0];
  assign reg_559__clk = clk;
  assign out_559[15:0] = reg_559__out[15:0];
  assign reg_56__clk = clk;
  assign out_56[15:0] = reg_56__out[15:0];
  assign reg_560__clk = clk;
  assign out_560[15:0] = reg_560__out[15:0];
  assign reg_561__clk = clk;
  assign out_561[15:0] = reg_561__out[15:0];
  assign reg_562__clk = clk;
  assign out_562[15:0] = reg_562__out[15:0];
  assign reg_563__clk = clk;
  assign out_563[15:0] = reg_563__out[15:0];
  assign reg_564__clk = clk;
  assign out_564[15:0] = reg_564__out[15:0];
  assign reg_565__clk = clk;
  assign out_565[15:0] = reg_565__out[15:0];
  assign reg_566__clk = clk;
  assign out_566[15:0] = reg_566__out[15:0];
  assign reg_567__clk = clk;
  assign out_567[15:0] = reg_567__out[15:0];
  assign reg_568__clk = clk;
  assign out_568[15:0] = reg_568__out[15:0];
  assign reg_569__clk = clk;
  assign out_569[15:0] = reg_569__out[15:0];
  assign reg_57__clk = clk;
  assign out_57[15:0] = reg_57__out[15:0];
  assign reg_570__clk = clk;
  assign out_570[15:0] = reg_570__out[15:0];
  assign reg_571__clk = clk;
  assign out_571[15:0] = reg_571__out[15:0];
  assign reg_572__clk = clk;
  assign out_572[15:0] = reg_572__out[15:0];
  assign reg_573__clk = clk;
  assign out_573[15:0] = reg_573__out[15:0];
  assign reg_574__clk = clk;
  assign out_574[15:0] = reg_574__out[15:0];
  assign reg_575__clk = clk;
  assign out_575[15:0] = reg_575__out[15:0];
  assign reg_576__clk = clk;
  assign out_576[15:0] = reg_576__out[15:0];
  assign reg_577__clk = clk;
  assign out_577[15:0] = reg_577__out[15:0];
  assign reg_578__clk = clk;
  assign out_578[15:0] = reg_578__out[15:0];
  assign reg_579__clk = clk;
  assign out_579[15:0] = reg_579__out[15:0];
  assign reg_58__clk = clk;
  assign out_58[15:0] = reg_58__out[15:0];
  assign reg_580__clk = clk;
  assign out_580[15:0] = reg_580__out[15:0];
  assign reg_581__clk = clk;
  assign out_581[15:0] = reg_581__out[15:0];
  assign reg_582__clk = clk;
  assign out_582[15:0] = reg_582__out[15:0];
  assign reg_583__clk = clk;
  assign out_583[15:0] = reg_583__out[15:0];
  assign reg_584__clk = clk;
  assign out_584[15:0] = reg_584__out[15:0];
  assign reg_585__clk = clk;
  assign out_585[15:0] = reg_585__out[15:0];
  assign reg_586__clk = clk;
  assign out_586[15:0] = reg_586__out[15:0];
  assign reg_587__clk = clk;
  assign out_587[15:0] = reg_587__out[15:0];
  assign reg_588__clk = clk;
  assign out_588[15:0] = reg_588__out[15:0];
  assign reg_589__clk = clk;
  assign out_589[15:0] = reg_589__out[15:0];
  assign reg_59__clk = clk;
  assign out_59[15:0] = reg_59__out[15:0];
  assign reg_590__clk = clk;
  assign out_590[15:0] = reg_590__out[15:0];
  assign reg_591__clk = clk;
  assign out_591[15:0] = reg_591__out[15:0];
  assign reg_592__clk = clk;
  assign out_592[15:0] = reg_592__out[15:0];
  assign reg_593__clk = clk;
  assign out_593[15:0] = reg_593__out[15:0];
  assign reg_594__clk = clk;
  assign out_594[15:0] = reg_594__out[15:0];
  assign reg_595__clk = clk;
  assign out_595[15:0] = reg_595__out[15:0];
  assign reg_596__clk = clk;
  assign out_596[15:0] = reg_596__out[15:0];
  assign reg_597__clk = clk;
  assign out_597[15:0] = reg_597__out[15:0];
  assign reg_598__clk = clk;
  assign out_598[15:0] = reg_598__out[15:0];
  assign reg_599__clk = clk;
  assign out_599[15:0] = reg_599__out[15:0];
  assign reg_6__clk = clk;
  assign out_6[15:0] = reg_6__out[15:0];
  assign reg_60__clk = clk;
  assign out_60[15:0] = reg_60__out[15:0];
  assign reg_600__clk = clk;
  assign out_600[15:0] = reg_600__out[15:0];
  assign reg_601__clk = clk;
  assign out_601[15:0] = reg_601__out[15:0];
  assign reg_602__clk = clk;
  assign out_602[15:0] = reg_602__out[15:0];
  assign reg_603__clk = clk;
  assign out_603[15:0] = reg_603__out[15:0];
  assign reg_604__clk = clk;
  assign out_604[15:0] = reg_604__out[15:0];
  assign reg_605__clk = clk;
  assign out_605[15:0] = reg_605__out[15:0];
  assign reg_606__clk = clk;
  assign out_606[15:0] = reg_606__out[15:0];
  assign reg_607__clk = clk;
  assign out_607[15:0] = reg_607__out[15:0];
  assign reg_608__clk = clk;
  assign out_608[15:0] = reg_608__out[15:0];
  assign reg_609__clk = clk;
  assign out_609[15:0] = reg_609__out[15:0];
  assign reg_61__clk = clk;
  assign out_61[15:0] = reg_61__out[15:0];
  assign reg_610__clk = clk;
  assign out_610[15:0] = reg_610__out[15:0];
  assign reg_611__clk = clk;
  assign out_611[15:0] = reg_611__out[15:0];
  assign reg_612__clk = clk;
  assign out_612[15:0] = reg_612__out[15:0];
  assign reg_613__clk = clk;
  assign out_613[15:0] = reg_613__out[15:0];
  assign reg_614__clk = clk;
  assign out_614[15:0] = reg_614__out[15:0];
  assign reg_615__clk = clk;
  assign out_615[15:0] = reg_615__out[15:0];
  assign reg_616__clk = clk;
  assign out_616[15:0] = reg_616__out[15:0];
  assign reg_617__clk = clk;
  assign out_617[15:0] = reg_617__out[15:0];
  assign reg_618__clk = clk;
  assign out_618[15:0] = reg_618__out[15:0];
  assign reg_619__clk = clk;
  assign out_619[15:0] = reg_619__out[15:0];
  assign reg_62__clk = clk;
  assign out_62[15:0] = reg_62__out[15:0];
  assign reg_620__clk = clk;
  assign out_620[15:0] = reg_620__out[15:0];
  assign reg_621__clk = clk;
  assign out_621[15:0] = reg_621__out[15:0];
  assign reg_622__clk = clk;
  assign out_622[15:0] = reg_622__out[15:0];
  assign reg_623__clk = clk;
  assign out_623[15:0] = reg_623__out[15:0];
  assign reg_624__clk = clk;
  assign out_624[15:0] = reg_624__out[15:0];
  assign reg_625__clk = clk;
  assign out_625[15:0] = reg_625__out[15:0];
  assign reg_626__clk = clk;
  assign out_626[15:0] = reg_626__out[15:0];
  assign reg_627__clk = clk;
  assign out_627[15:0] = reg_627__out[15:0];
  assign reg_628__clk = clk;
  assign out_628[15:0] = reg_628__out[15:0];
  assign reg_629__clk = clk;
  assign out_629[15:0] = reg_629__out[15:0];
  assign reg_63__clk = clk;
  assign out_63[15:0] = reg_63__out[15:0];
  assign reg_630__clk = clk;
  assign out_630[15:0] = reg_630__out[15:0];
  assign reg_631__clk = clk;
  assign out_631[15:0] = reg_631__out[15:0];
  assign reg_632__clk = clk;
  assign out_632[15:0] = reg_632__out[15:0];
  assign reg_633__clk = clk;
  assign out_633[15:0] = reg_633__out[15:0];
  assign reg_634__clk = clk;
  assign out_634[15:0] = reg_634__out[15:0];
  assign reg_635__clk = clk;
  assign out_635[15:0] = reg_635__out[15:0];
  assign reg_636__clk = clk;
  assign out_636[15:0] = reg_636__out[15:0];
  assign reg_637__clk = clk;
  assign out_637[15:0] = reg_637__out[15:0];
  assign reg_638__clk = clk;
  assign out_638[15:0] = reg_638__out[15:0];
  assign reg_639__clk = clk;
  assign out_639[15:0] = reg_639__out[15:0];
  assign reg_64__clk = clk;
  assign out_64[15:0] = reg_64__out[15:0];
  assign reg_640__clk = clk;
  assign out_640[15:0] = reg_640__out[15:0];
  assign reg_641__clk = clk;
  assign out_641[15:0] = reg_641__out[15:0];
  assign reg_642__clk = clk;
  assign out_642[15:0] = reg_642__out[15:0];
  assign reg_643__clk = clk;
  assign out_643[15:0] = reg_643__out[15:0];
  assign reg_644__clk = clk;
  assign out_644[15:0] = reg_644__out[15:0];
  assign reg_645__clk = clk;
  assign out_645[15:0] = reg_645__out[15:0];
  assign reg_646__clk = clk;
  assign out_646[15:0] = reg_646__out[15:0];
  assign reg_647__clk = clk;
  assign out_647[15:0] = reg_647__out[15:0];
  assign reg_648__clk = clk;
  assign out_648[15:0] = reg_648__out[15:0];
  assign reg_649__clk = clk;
  assign out_649[15:0] = reg_649__out[15:0];
  assign reg_65__clk = clk;
  assign out_65[15:0] = reg_65__out[15:0];
  assign reg_650__clk = clk;
  assign out_650[15:0] = reg_650__out[15:0];
  assign reg_651__clk = clk;
  assign out_651[15:0] = reg_651__out[15:0];
  assign reg_652__clk = clk;
  assign out_652[15:0] = reg_652__out[15:0];
  assign reg_653__clk = clk;
  assign out_653[15:0] = reg_653__out[15:0];
  assign reg_654__clk = clk;
  assign out_654[15:0] = reg_654__out[15:0];
  assign reg_655__clk = clk;
  assign out_655[15:0] = reg_655__out[15:0];
  assign reg_656__clk = clk;
  assign out_656[15:0] = reg_656__out[15:0];
  assign reg_657__clk = clk;
  assign out_657[15:0] = reg_657__out[15:0];
  assign reg_658__clk = clk;
  assign out_658[15:0] = reg_658__out[15:0];
  assign reg_659__clk = clk;
  assign out_659[15:0] = reg_659__out[15:0];
  assign reg_66__clk = clk;
  assign out_66[15:0] = reg_66__out[15:0];
  assign reg_660__clk = clk;
  assign out_660[15:0] = reg_660__out[15:0];
  assign reg_661__clk = clk;
  assign out_661[15:0] = reg_661__out[15:0];
  assign reg_662__clk = clk;
  assign out_662[15:0] = reg_662__out[15:0];
  assign reg_663__clk = clk;
  assign out_663[15:0] = reg_663__out[15:0];
  assign reg_664__clk = clk;
  assign out_664[15:0] = reg_664__out[15:0];
  assign reg_665__clk = clk;
  assign out_665[15:0] = reg_665__out[15:0];
  assign reg_666__clk = clk;
  assign out_666[15:0] = reg_666__out[15:0];
  assign reg_667__clk = clk;
  assign out_667[15:0] = reg_667__out[15:0];
  assign reg_668__clk = clk;
  assign out_668[15:0] = reg_668__out[15:0];
  assign reg_669__clk = clk;
  assign out_669[15:0] = reg_669__out[15:0];
  assign reg_67__clk = clk;
  assign out_67[15:0] = reg_67__out[15:0];
  assign reg_670__clk = clk;
  assign out_670[15:0] = reg_670__out[15:0];
  assign reg_671__clk = clk;
  assign out_671[15:0] = reg_671__out[15:0];
  assign reg_672__clk = clk;
  assign out_672[15:0] = reg_672__out[15:0];
  assign reg_673__clk = clk;
  assign out_673[15:0] = reg_673__out[15:0];
  assign reg_674__clk = clk;
  assign out_674[15:0] = reg_674__out[15:0];
  assign reg_675__clk = clk;
  assign out_675[15:0] = reg_675__out[15:0];
  assign reg_676__clk = clk;
  assign out_676[15:0] = reg_676__out[15:0];
  assign reg_677__clk = clk;
  assign out_677[15:0] = reg_677__out[15:0];
  assign reg_678__clk = clk;
  assign out_678[15:0] = reg_678__out[15:0];
  assign reg_679__clk = clk;
  assign out_679[15:0] = reg_679__out[15:0];
  assign reg_68__clk = clk;
  assign out_68[15:0] = reg_68__out[15:0];
  assign reg_680__clk = clk;
  assign out_680[15:0] = reg_680__out[15:0];
  assign reg_681__clk = clk;
  assign out_681[15:0] = reg_681__out[15:0];
  assign reg_682__clk = clk;
  assign out_682[15:0] = reg_682__out[15:0];
  assign reg_683__clk = clk;
  assign out_683[15:0] = reg_683__out[15:0];
  assign reg_684__clk = clk;
  assign out_684[15:0] = reg_684__out[15:0];
  assign reg_685__clk = clk;
  assign out_685[15:0] = reg_685__out[15:0];
  assign reg_686__clk = clk;
  assign out_686[15:0] = reg_686__out[15:0];
  assign reg_687__clk = clk;
  assign out_687[15:0] = reg_687__out[15:0];
  assign reg_688__clk = clk;
  assign out_688[15:0] = reg_688__out[15:0];
  assign reg_689__clk = clk;
  assign out_689[15:0] = reg_689__out[15:0];
  assign reg_69__clk = clk;
  assign out_69[15:0] = reg_69__out[15:0];
  assign reg_690__clk = clk;
  assign out_690[15:0] = reg_690__out[15:0];
  assign reg_691__clk = clk;
  assign out_691[15:0] = reg_691__out[15:0];
  assign reg_692__clk = clk;
  assign out_692[15:0] = reg_692__out[15:0];
  assign reg_693__clk = clk;
  assign out_693[15:0] = reg_693__out[15:0];
  assign reg_694__clk = clk;
  assign out_694[15:0] = reg_694__out[15:0];
  assign reg_695__clk = clk;
  assign out_695[15:0] = reg_695__out[15:0];
  assign reg_696__clk = clk;
  assign out_696[15:0] = reg_696__out[15:0];
  assign reg_697__clk = clk;
  assign out_697[15:0] = reg_697__out[15:0];
  assign reg_698__clk = clk;
  assign out_698[15:0] = reg_698__out[15:0];
  assign reg_699__clk = clk;
  assign out_699[15:0] = reg_699__out[15:0];
  assign reg_7__clk = clk;
  assign out_7[15:0] = reg_7__out[15:0];
  assign reg_70__clk = clk;
  assign out_70[15:0] = reg_70__out[15:0];
  assign reg_700__clk = clk;
  assign out_700[15:0] = reg_700__out[15:0];
  assign reg_701__clk = clk;
  assign out_701[15:0] = reg_701__out[15:0];
  assign reg_702__clk = clk;
  assign out_702[15:0] = reg_702__out[15:0];
  assign reg_703__clk = clk;
  assign out_703[15:0] = reg_703__out[15:0];
  assign reg_704__clk = clk;
  assign out_704[15:0] = reg_704__out[15:0];
  assign reg_705__clk = clk;
  assign out_705[15:0] = reg_705__out[15:0];
  assign reg_706__clk = clk;
  assign out_706[15:0] = reg_706__out[15:0];
  assign reg_707__clk = clk;
  assign out_707[15:0] = reg_707__out[15:0];
  assign reg_708__clk = clk;
  assign out_708[15:0] = reg_708__out[15:0];
  assign reg_709__clk = clk;
  assign out_709[15:0] = reg_709__out[15:0];
  assign reg_71__clk = clk;
  assign out_71[15:0] = reg_71__out[15:0];
  assign reg_710__clk = clk;
  assign out_710[15:0] = reg_710__out[15:0];
  assign reg_711__clk = clk;
  assign out_711[15:0] = reg_711__out[15:0];
  assign reg_712__clk = clk;
  assign out_712[15:0] = reg_712__out[15:0];
  assign reg_713__clk = clk;
  assign out_713[15:0] = reg_713__out[15:0];
  assign reg_714__clk = clk;
  assign out_714[15:0] = reg_714__out[15:0];
  assign reg_715__clk = clk;
  assign out_715[15:0] = reg_715__out[15:0];
  assign reg_716__clk = clk;
  assign out_716[15:0] = reg_716__out[15:0];
  assign reg_717__clk = clk;
  assign out_717[15:0] = reg_717__out[15:0];
  assign reg_718__clk = clk;
  assign out_718[15:0] = reg_718__out[15:0];
  assign reg_719__clk = clk;
  assign out_719[15:0] = reg_719__out[15:0];
  assign reg_72__clk = clk;
  assign out_72[15:0] = reg_72__out[15:0];
  assign reg_720__clk = clk;
  assign out_720[15:0] = reg_720__out[15:0];
  assign reg_721__clk = clk;
  assign out_721[15:0] = reg_721__out[15:0];
  assign reg_722__clk = clk;
  assign out_722[15:0] = reg_722__out[15:0];
  assign reg_723__clk = clk;
  assign out_723[15:0] = reg_723__out[15:0];
  assign reg_724__clk = clk;
  assign out_724[15:0] = reg_724__out[15:0];
  assign reg_725__clk = clk;
  assign out_725[15:0] = reg_725__out[15:0];
  assign reg_726__clk = clk;
  assign out_726[15:0] = reg_726__out[15:0];
  assign reg_727__clk = clk;
  assign out_727[15:0] = reg_727__out[15:0];
  assign reg_728__clk = clk;
  assign out_728[15:0] = reg_728__out[15:0];
  assign reg_729__clk = clk;
  assign out_729[15:0] = reg_729__out[15:0];
  assign reg_73__clk = clk;
  assign out_73[15:0] = reg_73__out[15:0];
  assign reg_730__clk = clk;
  assign out_730[15:0] = reg_730__out[15:0];
  assign reg_731__clk = clk;
  assign out_731[15:0] = reg_731__out[15:0];
  assign reg_732__clk = clk;
  assign out_732[15:0] = reg_732__out[15:0];
  assign reg_733__clk = clk;
  assign out_733[15:0] = reg_733__out[15:0];
  assign reg_734__clk = clk;
  assign out_734[15:0] = reg_734__out[15:0];
  assign reg_735__clk = clk;
  assign out_735[15:0] = reg_735__out[15:0];
  assign reg_736__clk = clk;
  assign out_736[15:0] = reg_736__out[15:0];
  assign reg_737__clk = clk;
  assign out_737[15:0] = reg_737__out[15:0];
  assign reg_738__clk = clk;
  assign out_738[15:0] = reg_738__out[15:0];
  assign reg_739__clk = clk;
  assign out_739[15:0] = reg_739__out[15:0];
  assign reg_74__clk = clk;
  assign out_74[15:0] = reg_74__out[15:0];
  assign reg_740__clk = clk;
  assign out_740[15:0] = reg_740__out[15:0];
  assign reg_741__clk = clk;
  assign out_741[15:0] = reg_741__out[15:0];
  assign reg_742__clk = clk;
  assign out_742[15:0] = reg_742__out[15:0];
  assign reg_743__clk = clk;
  assign out_743[15:0] = reg_743__out[15:0];
  assign reg_744__clk = clk;
  assign out_744[15:0] = reg_744__out[15:0];
  assign reg_745__clk = clk;
  assign out_745[15:0] = reg_745__out[15:0];
  assign reg_746__clk = clk;
  assign out_746[15:0] = reg_746__out[15:0];
  assign reg_747__clk = clk;
  assign out_747[15:0] = reg_747__out[15:0];
  assign reg_748__clk = clk;
  assign out_748[15:0] = reg_748__out[15:0];
  assign reg_749__clk = clk;
  assign out_749[15:0] = reg_749__out[15:0];
  assign reg_75__clk = clk;
  assign out_75[15:0] = reg_75__out[15:0];
  assign reg_750__clk = clk;
  assign out_750[15:0] = reg_750__out[15:0];
  assign reg_751__clk = clk;
  assign out_751[15:0] = reg_751__out[15:0];
  assign reg_752__clk = clk;
  assign out_752[15:0] = reg_752__out[15:0];
  assign reg_753__clk = clk;
  assign out_753[15:0] = reg_753__out[15:0];
  assign reg_754__clk = clk;
  assign out_754[15:0] = reg_754__out[15:0];
  assign reg_755__clk = clk;
  assign out_755[15:0] = reg_755__out[15:0];
  assign reg_756__clk = clk;
  assign out_756[15:0] = reg_756__out[15:0];
  assign reg_757__clk = clk;
  assign out_757[15:0] = reg_757__out[15:0];
  assign reg_758__clk = clk;
  assign out_758[15:0] = reg_758__out[15:0];
  assign reg_759__clk = clk;
  assign out_759[15:0] = reg_759__out[15:0];
  assign reg_76__clk = clk;
  assign out_76[15:0] = reg_76__out[15:0];
  assign reg_760__clk = clk;
  assign out_760[15:0] = reg_760__out[15:0];
  assign reg_761__clk = clk;
  assign out_761[15:0] = reg_761__out[15:0];
  assign reg_762__clk = clk;
  assign out_762[15:0] = reg_762__out[15:0];
  assign reg_763__clk = clk;
  assign out_763[15:0] = reg_763__out[15:0];
  assign reg_764__clk = clk;
  assign out_764[15:0] = reg_764__out[15:0];
  assign reg_765__clk = clk;
  assign out_765[15:0] = reg_765__out[15:0];
  assign reg_766__clk = clk;
  assign out_766[15:0] = reg_766__out[15:0];
  assign reg_767__clk = clk;
  assign out_767[15:0] = reg_767__out[15:0];
  assign reg_768__clk = clk;
  assign out_768[15:0] = reg_768__out[15:0];
  assign reg_769__clk = clk;
  assign out_769[15:0] = reg_769__out[15:0];
  assign reg_77__clk = clk;
  assign out_77[15:0] = reg_77__out[15:0];
  assign reg_770__clk = clk;
  assign out_770[15:0] = reg_770__out[15:0];
  assign reg_771__clk = clk;
  assign out_771[15:0] = reg_771__out[15:0];
  assign reg_772__clk = clk;
  assign out_772[15:0] = reg_772__out[15:0];
  assign reg_773__clk = clk;
  assign out_773[15:0] = reg_773__out[15:0];
  assign reg_774__clk = clk;
  assign out_774[15:0] = reg_774__out[15:0];
  assign reg_775__clk = clk;
  assign out_775[15:0] = reg_775__out[15:0];
  assign reg_776__clk = clk;
  assign out_776[15:0] = reg_776__out[15:0];
  assign reg_777__clk = clk;
  assign out_777[15:0] = reg_777__out[15:0];
  assign reg_778__clk = clk;
  assign out_778[15:0] = reg_778__out[15:0];
  assign reg_779__clk = clk;
  assign out_779[15:0] = reg_779__out[15:0];
  assign reg_78__clk = clk;
  assign out_78[15:0] = reg_78__out[15:0];
  assign reg_780__clk = clk;
  assign out_780[15:0] = reg_780__out[15:0];
  assign reg_781__clk = clk;
  assign out_781[15:0] = reg_781__out[15:0];
  assign reg_782__clk = clk;
  assign out_782[15:0] = reg_782__out[15:0];
  assign reg_783__clk = clk;
  assign out_783[15:0] = reg_783__out[15:0];
  assign reg_784__clk = clk;
  assign out_784[15:0] = reg_784__out[15:0];
  assign reg_785__clk = clk;
  assign out_785[15:0] = reg_785__out[15:0];
  assign reg_786__clk = clk;
  assign out_786[15:0] = reg_786__out[15:0];
  assign reg_787__clk = clk;
  assign out_787[15:0] = reg_787__out[15:0];
  assign reg_788__clk = clk;
  assign out_788[15:0] = reg_788__out[15:0];
  assign reg_789__clk = clk;
  assign out_789[15:0] = reg_789__out[15:0];
  assign reg_79__clk = clk;
  assign out_79[15:0] = reg_79__out[15:0];
  assign reg_790__clk = clk;
  assign out_790[15:0] = reg_790__out[15:0];
  assign reg_791__clk = clk;
  assign out_791[15:0] = reg_791__out[15:0];
  assign reg_792__clk = clk;
  assign out_792[15:0] = reg_792__out[15:0];
  assign reg_793__clk = clk;
  assign out_793[15:0] = reg_793__out[15:0];
  assign reg_794__clk = clk;
  assign out_794[15:0] = reg_794__out[15:0];
  assign reg_795__clk = clk;
  assign out_795[15:0] = reg_795__out[15:0];
  assign reg_796__clk = clk;
  assign out_796[15:0] = reg_796__out[15:0];
  assign reg_797__clk = clk;
  assign out_797[15:0] = reg_797__out[15:0];
  assign reg_798__clk = clk;
  assign out_798[15:0] = reg_798__out[15:0];
  assign reg_799__clk = clk;
  assign out_799[15:0] = reg_799__out[15:0];
  assign reg_8__clk = clk;
  assign out_8[15:0] = reg_8__out[15:0];
  assign reg_80__clk = clk;
  assign out_80[15:0] = reg_80__out[15:0];
  assign reg_800__clk = clk;
  assign out_800[15:0] = reg_800__out[15:0];
  assign reg_801__clk = clk;
  assign out_801[15:0] = reg_801__out[15:0];
  assign reg_802__clk = clk;
  assign out_802[15:0] = reg_802__out[15:0];
  assign reg_803__clk = clk;
  assign out_803[15:0] = reg_803__out[15:0];
  assign reg_804__clk = clk;
  assign out_804[15:0] = reg_804__out[15:0];
  assign reg_805__clk = clk;
  assign out_805[15:0] = reg_805__out[15:0];
  assign reg_806__clk = clk;
  assign out_806[15:0] = reg_806__out[15:0];
  assign reg_807__clk = clk;
  assign out_807[15:0] = reg_807__out[15:0];
  assign reg_808__clk = clk;
  assign out_808[15:0] = reg_808__out[15:0];
  assign reg_809__clk = clk;
  assign out_809[15:0] = reg_809__out[15:0];
  assign reg_81__clk = clk;
  assign out_81[15:0] = reg_81__out[15:0];
  assign reg_810__clk = clk;
  assign out_810[15:0] = reg_810__out[15:0];
  assign reg_811__clk = clk;
  assign out_811[15:0] = reg_811__out[15:0];
  assign reg_812__clk = clk;
  assign out_812[15:0] = reg_812__out[15:0];
  assign reg_813__clk = clk;
  assign out_813[15:0] = reg_813__out[15:0];
  assign reg_814__clk = clk;
  assign out_814[15:0] = reg_814__out[15:0];
  assign reg_815__clk = clk;
  assign out_815[15:0] = reg_815__out[15:0];
  assign reg_816__clk = clk;
  assign out_816[15:0] = reg_816__out[15:0];
  assign reg_817__clk = clk;
  assign out_817[15:0] = reg_817__out[15:0];
  assign reg_818__clk = clk;
  assign out_818[15:0] = reg_818__out[15:0];
  assign reg_819__clk = clk;
  assign out_819[15:0] = reg_819__out[15:0];
  assign reg_82__clk = clk;
  assign out_82[15:0] = reg_82__out[15:0];
  assign reg_820__clk = clk;
  assign out_820[15:0] = reg_820__out[15:0];
  assign reg_821__clk = clk;
  assign out_821[15:0] = reg_821__out[15:0];
  assign reg_822__clk = clk;
  assign out_822[15:0] = reg_822__out[15:0];
  assign reg_823__clk = clk;
  assign out_823[15:0] = reg_823__out[15:0];
  assign reg_824__clk = clk;
  assign out_824[15:0] = reg_824__out[15:0];
  assign reg_825__clk = clk;
  assign out_825[15:0] = reg_825__out[15:0];
  assign reg_826__clk = clk;
  assign out_826[15:0] = reg_826__out[15:0];
  assign reg_827__clk = clk;
  assign out_827[15:0] = reg_827__out[15:0];
  assign reg_828__clk = clk;
  assign out_828[15:0] = reg_828__out[15:0];
  assign reg_829__clk = clk;
  assign out_829[15:0] = reg_829__out[15:0];
  assign reg_83__clk = clk;
  assign out_83[15:0] = reg_83__out[15:0];
  assign reg_830__clk = clk;
  assign out_830[15:0] = reg_830__out[15:0];
  assign reg_831__clk = clk;
  assign out_831[15:0] = reg_831__out[15:0];
  assign reg_832__clk = clk;
  assign out_832[15:0] = reg_832__out[15:0];
  assign reg_833__clk = clk;
  assign out_833[15:0] = reg_833__out[15:0];
  assign reg_834__clk = clk;
  assign out_834[15:0] = reg_834__out[15:0];
  assign reg_835__clk = clk;
  assign out_835[15:0] = reg_835__out[15:0];
  assign reg_836__clk = clk;
  assign out_836[15:0] = reg_836__out[15:0];
  assign reg_837__clk = clk;
  assign out_837[15:0] = reg_837__out[15:0];
  assign reg_838__clk = clk;
  assign out_838[15:0] = reg_838__out[15:0];
  assign reg_839__clk = clk;
  assign out_839[15:0] = reg_839__out[15:0];
  assign reg_84__clk = clk;
  assign out_84[15:0] = reg_84__out[15:0];
  assign reg_840__clk = clk;
  assign out_840[15:0] = reg_840__out[15:0];
  assign reg_841__clk = clk;
  assign out_841[15:0] = reg_841__out[15:0];
  assign reg_842__clk = clk;
  assign out_842[15:0] = reg_842__out[15:0];
  assign reg_843__clk = clk;
  assign out_843[15:0] = reg_843__out[15:0];
  assign reg_844__clk = clk;
  assign out_844[15:0] = reg_844__out[15:0];
  assign reg_845__clk = clk;
  assign out_845[15:0] = reg_845__out[15:0];
  assign reg_846__clk = clk;
  assign out_846[15:0] = reg_846__out[15:0];
  assign reg_847__clk = clk;
  assign out_847[15:0] = reg_847__out[15:0];
  assign reg_848__clk = clk;
  assign out_848[15:0] = reg_848__out[15:0];
  assign reg_849__clk = clk;
  assign out_849[15:0] = reg_849__out[15:0];
  assign reg_85__clk = clk;
  assign out_85[15:0] = reg_85__out[15:0];
  assign reg_850__clk = clk;
  assign out_850[15:0] = reg_850__out[15:0];
  assign reg_851__clk = clk;
  assign out_851[15:0] = reg_851__out[15:0];
  assign reg_852__clk = clk;
  assign out_852[15:0] = reg_852__out[15:0];
  assign reg_853__clk = clk;
  assign out_853[15:0] = reg_853__out[15:0];
  assign reg_854__clk = clk;
  assign out_854[15:0] = reg_854__out[15:0];
  assign reg_855__clk = clk;
  assign out_855[15:0] = reg_855__out[15:0];
  assign reg_856__clk = clk;
  assign out_856[15:0] = reg_856__out[15:0];
  assign reg_857__clk = clk;
  assign out_857[15:0] = reg_857__out[15:0];
  assign reg_858__clk = clk;
  assign out_858[15:0] = reg_858__out[15:0];
  assign reg_859__clk = clk;
  assign out_859[15:0] = reg_859__out[15:0];
  assign reg_86__clk = clk;
  assign out_86[15:0] = reg_86__out[15:0];
  assign reg_860__clk = clk;
  assign out_860[15:0] = reg_860__out[15:0];
  assign reg_861__clk = clk;
  assign out_861[15:0] = reg_861__out[15:0];
  assign reg_862__clk = clk;
  assign out_862[15:0] = reg_862__out[15:0];
  assign reg_863__clk = clk;
  assign out_863[15:0] = reg_863__out[15:0];
  assign reg_864__clk = clk;
  assign out_864[15:0] = reg_864__out[15:0];
  assign reg_865__clk = clk;
  assign out_865[15:0] = reg_865__out[15:0];
  assign reg_866__clk = clk;
  assign out_866[15:0] = reg_866__out[15:0];
  assign reg_867__clk = clk;
  assign out_867[15:0] = reg_867__out[15:0];
  assign reg_868__clk = clk;
  assign out_868[15:0] = reg_868__out[15:0];
  assign reg_869__clk = clk;
  assign out_869[15:0] = reg_869__out[15:0];
  assign reg_87__clk = clk;
  assign out_87[15:0] = reg_87__out[15:0];
  assign reg_870__clk = clk;
  assign out_870[15:0] = reg_870__out[15:0];
  assign reg_871__clk = clk;
  assign out_871[15:0] = reg_871__out[15:0];
  assign reg_872__clk = clk;
  assign out_872[15:0] = reg_872__out[15:0];
  assign reg_873__clk = clk;
  assign out_873[15:0] = reg_873__out[15:0];
  assign reg_874__clk = clk;
  assign out_874[15:0] = reg_874__out[15:0];
  assign reg_875__clk = clk;
  assign out_875[15:0] = reg_875__out[15:0];
  assign reg_876__clk = clk;
  assign out_876[15:0] = reg_876__out[15:0];
  assign reg_877__clk = clk;
  assign out_877[15:0] = reg_877__out[15:0];
  assign reg_878__clk = clk;
  assign out_878[15:0] = reg_878__out[15:0];
  assign reg_879__clk = clk;
  assign out_879[15:0] = reg_879__out[15:0];
  assign reg_88__clk = clk;
  assign out_88[15:0] = reg_88__out[15:0];
  assign reg_880__clk = clk;
  assign out_880[15:0] = reg_880__out[15:0];
  assign reg_881__clk = clk;
  assign out_881[15:0] = reg_881__out[15:0];
  assign reg_882__clk = clk;
  assign out_882[15:0] = reg_882__out[15:0];
  assign reg_883__clk = clk;
  assign out_883[15:0] = reg_883__out[15:0];
  assign reg_884__clk = clk;
  assign out_884[15:0] = reg_884__out[15:0];
  assign reg_885__clk = clk;
  assign out_885[15:0] = reg_885__out[15:0];
  assign reg_886__clk = clk;
  assign out_886[15:0] = reg_886__out[15:0];
  assign reg_887__clk = clk;
  assign out_887[15:0] = reg_887__out[15:0];
  assign reg_888__clk = clk;
  assign out_888[15:0] = reg_888__out[15:0];
  assign reg_889__clk = clk;
  assign out_889[15:0] = reg_889__out[15:0];
  assign reg_89__clk = clk;
  assign out_89[15:0] = reg_89__out[15:0];
  assign reg_890__clk = clk;
  assign out_890[15:0] = reg_890__out[15:0];
  assign reg_891__clk = clk;
  assign out_891[15:0] = reg_891__out[15:0];
  assign reg_892__clk = clk;
  assign out_892[15:0] = reg_892__out[15:0];
  assign reg_893__clk = clk;
  assign out_893[15:0] = reg_893__out[15:0];
  assign reg_894__clk = clk;
  assign out_894[15:0] = reg_894__out[15:0];
  assign reg_895__clk = clk;
  assign out_895[15:0] = reg_895__out[15:0];
  assign reg_896__clk = clk;
  assign out_896[15:0] = reg_896__out[15:0];
  assign reg_897__clk = clk;
  assign out_897[15:0] = reg_897__out[15:0];
  assign reg_898__clk = clk;
  assign out_898[15:0] = reg_898__out[15:0];
  assign reg_899__clk = clk;
  assign out_899[15:0] = reg_899__out[15:0];
  assign reg_9__clk = clk;
  assign out_9[15:0] = reg_9__out[15:0];
  assign reg_90__clk = clk;
  assign out_90[15:0] = reg_90__out[15:0];
  assign reg_900__clk = clk;
  assign out_900[15:0] = reg_900__out[15:0];
  assign reg_901__clk = clk;
  assign out_901[15:0] = reg_901__out[15:0];
  assign reg_902__clk = clk;
  assign out_902[15:0] = reg_902__out[15:0];
  assign reg_903__clk = clk;
  assign out_903[15:0] = reg_903__out[15:0];
  assign reg_904__clk = clk;
  assign out_904[15:0] = reg_904__out[15:0];
  assign reg_905__clk = clk;
  assign out_905[15:0] = reg_905__out[15:0];
  assign reg_906__clk = clk;
  assign out_906[15:0] = reg_906__out[15:0];
  assign reg_907__clk = clk;
  assign out_907[15:0] = reg_907__out[15:0];
  assign reg_908__clk = clk;
  assign out_908[15:0] = reg_908__out[15:0];
  assign reg_909__clk = clk;
  assign out_909[15:0] = reg_909__out[15:0];
  assign reg_91__clk = clk;
  assign out_91[15:0] = reg_91__out[15:0];
  assign reg_910__clk = clk;
  assign out_910[15:0] = reg_910__out[15:0];
  assign reg_911__clk = clk;
  assign out_911[15:0] = reg_911__out[15:0];
  assign reg_912__clk = clk;
  assign out_912[15:0] = reg_912__out[15:0];
  assign reg_913__clk = clk;
  assign out_913[15:0] = reg_913__out[15:0];
  assign reg_914__clk = clk;
  assign out_914[15:0] = reg_914__out[15:0];
  assign reg_915__clk = clk;
  assign out_915[15:0] = reg_915__out[15:0];
  assign reg_916__clk = clk;
  assign out_916[15:0] = reg_916__out[15:0];
  assign reg_917__clk = clk;
  assign out_917[15:0] = reg_917__out[15:0];
  assign reg_918__clk = clk;
  assign out_918[15:0] = reg_918__out[15:0];
  assign reg_919__clk = clk;
  assign out_919[15:0] = reg_919__out[15:0];
  assign reg_92__clk = clk;
  assign out_92[15:0] = reg_92__out[15:0];
  assign reg_920__clk = clk;
  assign out_920[15:0] = reg_920__out[15:0];
  assign reg_921__clk = clk;
  assign out_921[15:0] = reg_921__out[15:0];
  assign reg_922__clk = clk;
  assign out_922[15:0] = reg_922__out[15:0];
  assign reg_923__clk = clk;
  assign out_923[15:0] = reg_923__out[15:0];
  assign reg_924__clk = clk;
  assign out_924[15:0] = reg_924__out[15:0];
  assign reg_925__clk = clk;
  assign out_925[15:0] = reg_925__out[15:0];
  assign reg_926__clk = clk;
  assign out_926[15:0] = reg_926__out[15:0];
  assign reg_927__clk = clk;
  assign out_927[15:0] = reg_927__out[15:0];
  assign reg_928__clk = clk;
  assign out_928[15:0] = reg_928__out[15:0];
  assign reg_929__clk = clk;
  assign out_929[15:0] = reg_929__out[15:0];
  assign reg_93__clk = clk;
  assign out_93[15:0] = reg_93__out[15:0];
  assign reg_930__clk = clk;
  assign out_930[15:0] = reg_930__out[15:0];
  assign reg_931__clk = clk;
  assign out_931[15:0] = reg_931__out[15:0];
  assign reg_932__clk = clk;
  assign out_932[15:0] = reg_932__out[15:0];
  assign reg_933__clk = clk;
  assign out_933[15:0] = reg_933__out[15:0];
  assign reg_934__clk = clk;
  assign out_934[15:0] = reg_934__out[15:0];
  assign reg_935__clk = clk;
  assign out_935[15:0] = reg_935__out[15:0];
  assign reg_936__clk = clk;
  assign out_936[15:0] = reg_936__out[15:0];
  assign reg_937__clk = clk;
  assign out_937[15:0] = reg_937__out[15:0];
  assign reg_938__clk = clk;
  assign out_938[15:0] = reg_938__out[15:0];
  assign reg_939__clk = clk;
  assign out_939[15:0] = reg_939__out[15:0];
  assign reg_94__clk = clk;
  assign out_94[15:0] = reg_94__out[15:0];
  assign reg_940__clk = clk;
  assign out_940[15:0] = reg_940__out[15:0];
  assign reg_941__clk = clk;
  assign out_941[15:0] = reg_941__out[15:0];
  assign reg_942__clk = clk;
  assign out_942[15:0] = reg_942__out[15:0];
  assign reg_943__clk = clk;
  assign out_943[15:0] = reg_943__out[15:0];
  assign reg_944__clk = clk;
  assign out_944[15:0] = reg_944__out[15:0];
  assign reg_945__clk = clk;
  assign out_945[15:0] = reg_945__out[15:0];
  assign reg_946__clk = clk;
  assign out_946[15:0] = reg_946__out[15:0];
  assign reg_947__clk = clk;
  assign out_947[15:0] = reg_947__out[15:0];
  assign reg_948__clk = clk;
  assign out_948[15:0] = reg_948__out[15:0];
  assign reg_949__clk = clk;
  assign out_949[15:0] = reg_949__out[15:0];
  assign reg_95__clk = clk;
  assign out_95[15:0] = reg_95__out[15:0];
  assign reg_950__clk = clk;
  assign out_950[15:0] = reg_950__out[15:0];
  assign reg_951__clk = clk;
  assign out_951[15:0] = reg_951__out[15:0];
  assign reg_952__clk = clk;
  assign out_952[15:0] = reg_952__out[15:0];
  assign reg_953__clk = clk;
  assign out_953[15:0] = reg_953__out[15:0];
  assign reg_954__clk = clk;
  assign out_954[15:0] = reg_954__out[15:0];
  assign reg_955__clk = clk;
  assign out_955[15:0] = reg_955__out[15:0];
  assign reg_956__clk = clk;
  assign out_956[15:0] = reg_956__out[15:0];
  assign reg_957__clk = clk;
  assign out_957[15:0] = reg_957__out[15:0];
  assign reg_958__clk = clk;
  assign out_958[15:0] = reg_958__out[15:0];
  assign reg_959__clk = clk;
  assign out_959[15:0] = reg_959__out[15:0];
  assign reg_96__clk = clk;
  assign out_96[15:0] = reg_96__out[15:0];
  assign reg_960__clk = clk;
  assign out_960[15:0] = reg_960__out[15:0];
  assign reg_961__clk = clk;
  assign out_961[15:0] = reg_961__out[15:0];
  assign reg_962__clk = clk;
  assign out_962[15:0] = reg_962__out[15:0];
  assign reg_963__clk = clk;
  assign out_963[15:0] = reg_963__out[15:0];
  assign reg_964__clk = clk;
  assign out_964[15:0] = reg_964__out[15:0];
  assign reg_965__clk = clk;
  assign out_965[15:0] = reg_965__out[15:0];
  assign reg_966__clk = clk;
  assign out_966[15:0] = reg_966__out[15:0];
  assign reg_967__clk = clk;
  assign out_967[15:0] = reg_967__out[15:0];
  assign reg_968__clk = clk;
  assign out_968[15:0] = reg_968__out[15:0];
  assign reg_969__clk = clk;
  assign out_969[15:0] = reg_969__out[15:0];
  assign reg_97__clk = clk;
  assign out_97[15:0] = reg_97__out[15:0];
  assign reg_970__clk = clk;
  assign out_970[15:0] = reg_970__out[15:0];
  assign reg_971__clk = clk;
  assign out_971[15:0] = reg_971__out[15:0];
  assign reg_972__clk = clk;
  assign out_972[15:0] = reg_972__out[15:0];
  assign reg_973__clk = clk;
  assign out_973[15:0] = reg_973__out[15:0];
  assign reg_974__clk = clk;
  assign out_974[15:0] = reg_974__out[15:0];
  assign reg_975__clk = clk;
  assign out_975[15:0] = reg_975__out[15:0];
  assign reg_976__clk = clk;
  assign out_976[15:0] = reg_976__out[15:0];
  assign reg_977__clk = clk;
  assign out_977[15:0] = reg_977__out[15:0];
  assign reg_978__clk = clk;
  assign out_978[15:0] = reg_978__out[15:0];
  assign reg_979__clk = clk;
  assign out_979[15:0] = reg_979__out[15:0];
  assign reg_98__clk = clk;
  assign out_98[15:0] = reg_98__out[15:0];
  assign reg_980__clk = clk;
  assign out_980[15:0] = reg_980__out[15:0];
  assign reg_981__clk = clk;
  assign out_981[15:0] = reg_981__out[15:0];
  assign reg_982__clk = clk;
  assign out_982[15:0] = reg_982__out[15:0];
  assign reg_983__clk = clk;
  assign out_983[15:0] = reg_983__out[15:0];
  assign reg_984__clk = clk;
  assign out_984[15:0] = reg_984__out[15:0];
  assign reg_985__clk = clk;
  assign out_985[15:0] = reg_985__out[15:0];
  assign reg_986__clk = clk;
  assign out_986[15:0] = reg_986__out[15:0];
  assign reg_987__clk = clk;
  assign out_987[15:0] = reg_987__out[15:0];
  assign reg_988__clk = clk;
  assign out_988[15:0] = reg_988__out[15:0];
  assign reg_989__clk = clk;
  assign out_989[15:0] = reg_989__out[15:0];
  assign reg_99__clk = clk;
  assign out_99[15:0] = reg_99__out[15:0];
  assign reg_990__clk = clk;
  assign out_990[15:0] = reg_990__out[15:0];
  assign reg_991__clk = clk;
  assign out_991[15:0] = reg_991__out[15:0];
  assign reg_992__clk = clk;
  assign out_992[15:0] = reg_992__out[15:0];
  assign reg_993__clk = clk;
  assign out_993[15:0] = reg_993__out[15:0];
  assign reg_994__clk = clk;
  assign out_994[15:0] = reg_994__out[15:0];
  assign reg_995__clk = clk;
  assign out_995[15:0] = reg_995__out[15:0];
  assign reg_996__clk = clk;
  assign out_996[15:0] = reg_996__out[15:0];
  assign reg_997__clk = clk;
  assign out_997[15:0] = reg_997__out[15:0];
  assign reg_998__clk = clk;
  assign out_998[15:0] = reg_998__out[15:0];
  assign reg_999__clk = clk;
  assign out_999[15:0] = reg_999__out[15:0];

endmodule //manyOps
